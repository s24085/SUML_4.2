���/     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.2.2�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak��ST_Slope�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh&hNhJ�
hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��h4�f8�����R�(KhQNNNJ����J����K t�b�C              �?�t�bhUh(�scalar���hPC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hK�
node_count�K�nodes�h*h-K ��h/��R�(KK煔h4�V56�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h�h4�i8�����R�(KhQNNNJ����J����K t�bK ��h�h�K��h�h�K��h�haK��h�haK ��h�h�K(��h�haK0��uK8KKt�b�B�2         �                    �?j8je3�?�           ��@       G                    �?�}�	���?           �y@       6                   �a@�n_Y�K�?e            �c@       -       	          ����?     ^�?P             `@       $                    �?�/���?B            �Y@                          �_@�{��?5            �T@                           �?�q�q��?!             H@                           �?�4F����?            �D@	                          �c@z�G�z�?             @
                          �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?      �?             B@                          Pf@�q�q�?             "@������������������������       �                     @������������������������       �                     @                          �[@�<ݚ�?             ;@������������������������       �                     @              
             �?����X�?             5@������������������������       �                     *@                          @^@      �?              @������������������������       �                     @������������������������       �                      @                           �I@؇���X�?             @������������������������       �                     @                           @M@�q�q�?             @������������������������       �                     �?������������������������       �                      @       #       
             �?�t����?             A@       "                    �?���Q��?             $@        !                    �I@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     8@%       ,                    @L@���N8�?             5@&       +                   ``@�S����?             3@'       (                   n@�IєX�?             1@������������������������       �                     *@)       *                   �Y@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @.       /       	             �?`2U0*��?             9@������������������������       �                     $@0       5                    �H@��S�ۿ?	             .@1       2       
             �?      �?             @������������������������       �                      @3       4                   `T@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@7       F                   �y@�>4և��?             <@8       A       	             �?PN��T'�?             ;@9       @                   �e@      �?              @:       ?                   �b@����X�?             @;       <                   �`@      �?             @������������������������       �                     �?=       >       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?B       E                    �?�}�+r��?             3@C       D       
             �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     @������������������������       �                     �?H       �                    �?     ��?�             p@I       J                   �U@ ?����?w            @h@������������������������       �                     �?K       |                   �b@ː����?v             h@L       [                   �[@<;n,��?m             f@M       N                   �Y@z�G�z�?             >@������������������������       �                     @O       Z                   �m@��+7��?             7@P       Q                   ph@և���X�?             ,@������������������������       �                     @R       S                   �Z@�q�q�?             "@������������������������       �                      @T       Y                    b@և���X�?             @U       X                    �I@z�G�z�?             @V       W       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     "@\       s       
             �?�c!�^�?]            @b@]       ^                   �i@5�wAd�?T            �`@������������������������       �                     H@_       j                   �[@���1j	�?6            �U@`       i                    @M@<���D�?            �@@a       d                   `[@8�Z$���?             :@b       c                   0j@���N8�?             5@������������������������       �                     �?������������������������       �                     4@e       f                    �?���Q��?             @������������������������       �                     �?g       h                   �k@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @k       r       	          ����?�O4R���?!            �J@l       q                    �?�����H�?             "@m       n                   pb@z�G�z�?             @������������������������       �                      @o       p                   `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     F@t       {                    c@r�q��?	             (@u       z                    �?�C��2(�?             &@v       y                   �Z@r�q��?             @w       x                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?}       �       
             �?��.k���?	             1@~                          pn@���Q��?             $@������������������������       �                      @�       �                    q@      �?              @������������������������       �                     @������������������������       �                      @�       �                   `k@����X�?             @������������������������       �                     �?�       �                    �P@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �R@0�z��?�?%             O@������������������������       �        $            �N@������������������������       �                     �?�       �                    _@"\�����?�             t@�       �                    @K@�q�q�?,            @Q@�       �                   c@������?             1@�       �                    �?؇���X�?             ,@������������������������       �        	             &@�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    ^@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?���B���?             J@�       �       
             �?8^s]e�?             =@�       �                    `@�θ�?             :@������������������������       �                     &@�       �       	          pff�?���Q��?
             .@�       �                    @z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	          @33�?�nkK�?
             7@������������������������       �                     �?������������������������       �        	             6@�       �       	          033�?:]���?�            �o@�       �                    �?�iZi�?�             l@�       �                    @���I/��?�            @h@�       �       	          ����?`���i��?y             f@�       �       
             �?@+K&:~�?e             c@�       �                   �q@�t����?             1@�       �                   `]@      �?             0@������������������������       �                      @�       �                   �b@؇���X�?
             ,@������������������������       �                      @������������������������       �                     (@������������������������       �                     �?�       �       	          ����?`��(�?X            �`@�       �                   �t@�T�~~4�?M            @]@�       �                   h@����X�?I             \@������������������������       �        G            @[@�       �                    d@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@�       �                    �?�q�q�?             8@������������������������       �                     "@�       �                   �\@��S���?             .@������������������������       �                     @�       �                    �K@���!pc�?
             &@������������������������       �                     @�       �                    �M@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?b�2�tk�?             2@�       �                    �M@��S���?
             .@�       �                   �h@�<ݚ�?             "@�       �                   `e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   �`@�4�����?             ?@������������������������       �                     @�       �                     I@���B���?             :@������������������������       �                     @�       �       
             �?���7�?
             6@�       �                    �?z�G�z�?             @������������������������       �                     @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     1@�       �                    �?����X�?             <@������������������������       �                     @�       �       
             �?r�q��?             8@������������������������       �                     �?�       �                   @a@�LQ�1	�?             7@������������������������       �                     �?�       �                    c@�C��2(�?             6@������������������������       �                     &@�       �       	             @"pc�
�?             &@������������������������       �                     �?�       �                   Pd@ףp=
�?             $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�t�b�values�h*h-K ��h/��R�(KK�KK��ha�Bp       Ps@     �z@      U@     �t@      N@      X@     �K@     @R@      K@     �H@     �H@     �@@      3@      =@      *@      <@      @      �?      �?      �?      �?                      �?      @              "@      ;@      @      @              @      @              @      5@              @      @      .@              *@      @       @      @                       @      @      �?      @               @      �?              �?       @              >@      @      @      @      @      @              @      @               @              8@              @      0@      @      0@      �?      0@              *@      �?      @      �?                      @       @               @              �?      8@              $@      �?      ,@      �?      @               @      �?      �?              �?      �?                      &@      @      7@      @      7@      @      @       @      @       @       @              �?       @      �?              �?       @                      @      �?              �?      2@      �?      &@              &@      �?                      @      �?              8@      m@      7@     `e@      �?              6@     `e@      *@     `d@      @      8@              @      @      1@      @       @              @      @      @       @              @      @      @      �?      �?      �?      �?                      �?      @                       @              "@      @     `a@      @      `@              H@      @     @T@      @      =@      @      6@      �?      4@      �?                      4@      @       @      �?               @       @               @       @                      @      �?      J@      �?       @      �?      @               @      �?       @      �?                       @              @              F@       @      $@      �?      $@      �?      @      �?      �?      �?                      �?              @              @      �?              "@       @      @      @       @               @      @              @       @              @       @              �?      @      �?      @                      �?      �?     �N@             �N@      �?              l@     @X@      7@      G@      *@      @      (@       @      &@              �?       @               @      �?              �?       @               @      �?              $@      E@      "@      4@      @      4@              &@      @      "@       @       @               @       @              @      �?      @                      �?      @              �?      6@      �?                      6@     @i@     �I@     @h@      ?@     �e@      5@     @d@      ,@      b@      @      (@      @      (@      @               @      (@       @               @      (@                      �?     �`@       @     �\@       @     �[@      �?     @[@               @      �?       @                      �?      @      �?      @                      �?      2@              1@      @      "@               @      @              @       @      @      @              @      @              @      @              &@      @       @      @       @      @       @      �?       @                      �?              @      @              @              5@      $@              @      5@      @              @      5@      �?      @      �?      @              �?      �?              �?      �?              1@               @      4@      @              @      4@      �?              @      4@      �?               @      4@              &@       @      "@      �?              �?      "@      �?      �?              �?      �?                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ/��hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKم�h��Bx/         �       
             �?4�5����?�           ��@       E                    �?P� �&�?           @y@                           �?l��\��?�             q@              
             �?�	j*D�?            �C@������������������������       �                     @                           �?���|���?            �@@                           @O@X�<ݚ�?             ;@       	                   �Z@�eP*L��?             6@������������������������       �                     @
                          �c@p�ݯ��?             3@                           b@     ��?             0@              	             �?      �?             (@                          �_@ףp=
�?             $@                          �p@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @                           �?�!��?�             m@������������������������       �                     F@                          �U@$Q�q�?y            �g@������������������������       �                     �?       D                   Pz@P��a4�?x            �g@       A                    �R@a��_�?w            `g@       $                   �g@p��D��?u             g@                           �?`����֜?,            �Q@������������������������       �                    �G@        #                    �?�nkK�?             7@!       "                    `@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     &@%       &                    Z@���^���?I            �\@������������������������       �                     8@'       <       	          ����?|)����?<            �V@(       1                   �\@X�;�^o�?!            �K@)       0                    @J@      �?             0@*       /                    b@؇���X�?             ,@+       .                    �?�q�q�?             @,       -       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @2       ;       	             �?$�q-�?            �C@3       4                   �i@���!pc�?             &@������������������������       �                     �?5       :                    �?z�G�z�?             $@6       7                    �?����X�?             @������������������������       �                     @8       9                     K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     <@=       @                    ]@������?             B@>       ?                   �m@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     <@B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?F       U                   0i@���e��?X            �`@G       H                    @G@�T|n�q�?            �E@������������������������       �                      @I       P       	          `ff@,���i�?            �D@J       O                    �?Pa�	�?            �@@K       N                   �b@      �?             @L       M       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     =@Q       R                    �?      �?              @������������������������       �                     �?S       T                   c@և���X�?             @������������������������       �                     @������������������������       �                     @V       ]                    �?dWp,���?=            @V@W       \                   �d@�C��2(�?             6@X       [                   �Z@���N8�?             5@Y       Z                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@������������������������       �                     �?^       {                   �`@�#}7��?.            �P@_       `                   �j@��
P��?            �A@������������������������       �                     @a       h                   �b@     ��?             @@b       g                     N@�����H�?             "@c       d                    @M@z�G�z�?             @������������������������       �                     @e       f                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @i       x                    �L@�û��|�?             7@j       s       	             @�����?             3@k       r       	             �?z�G�z�?	             .@l       q                    ]@�q�q�?             "@m       n                    �?      �?             @������������������������       �                      @o       p                   pf@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @t       w                    �?      �?             @u       v                   (p@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?y       z                    [@      �?             @������������������������       �                     �?������������������������       �                     @|       }                    @N@     ��?             @@������������������������       �                     4@~       �                    �?�q�q�?
             (@       �                   �b@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   pb@      �?             @������������������������       �                     @������������������������       �                     @�       �                   @E@`}�?��?�            �t@�       �                    �?P����?             C@�       �                    �K@��Q��?             4@�       �                    ]@      �?              @������������������������       �                      @�       �                   `\@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �c@r�q��?             (@�       �                    �?�C��2(�?             &@������������������������       �                     @�       �       	             �?      �?             @�       �                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     2@�       �                    �?�@i����?�            @r@�       �                    �?��|�	��?6            �V@������������������������       �                     .@�       �                    �?��=A��?/             S@�       �       	          ��� @��+7��?             7@�       �                   �f@�GN�z�?             6@������������������������       �        
             1@������������������������       �                     @������������������������       �                     �?�       �                   �X@Ȩ�I��?"            �J@������������������������       �                      @�       �       	          hff�?������?!            �I@�       �                    �?$�q-�?            �C@�       �                   �c@ȵHPS!�?             :@������������������������       �                     4@�       �                    �G@      �?             @�       �                   @b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@�       �                   @b@      �?             (@�       �                   �`@�����H�?             "@������������������������       �                     @�       �                    @J@z�G�z�?             @������������������������       �                     @�       �                   Pc@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �t@t�e�í�?z             i@�       �                   �g@�Q �?w            �h@�       �                    @�-j'�?v             h@�       �       	          ���@����?l             f@�       �                   c@@�E��@�?k            �e@�       �                    @L@p�|�i�?1             S@�       �                   @[@ ������?(            �O@�       �                    Z@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        &             M@�       �                   Hp@8�Z$���?	             *@������������������������       �                     @�       �                    �?����X�?             @�       �                   �p@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �        :            �X@������������������������       �                      @�       �                   Pp@     ��?
             0@�       �                   �d@8�Z$���?             *@�       �                    a@����X�?             @�       �                    �?      �?             @�       �                    c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �N@���Q��?             @������������������������       �                     @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       �t@     y@     �R@     �t@      8@      o@      (@      ;@              @      (@      5@      (@      .@      (@      $@              @      (@      @      "@      @      "@      @      "@      �?      @      �?              �?      @              @                       @              @      @                      @              @      (@     �k@              F@      (@      f@      �?              &@      f@      $@      f@      "@      f@      �?     @Q@             �G@      �?      6@      �?      &@      �?                      &@              &@       @     �Z@              8@       @     �T@      @      H@      @      (@       @      (@       @      @       @      �?              �?       @                      @               @       @              @      B@      @       @      �?               @       @       @      @              @       @      �?              �?       @                      @              <@      �?     �A@      �?      @              @      �?                      <@      �?      �?      �?                      �?      �?              I@     �T@      @      B@       @              @      B@      �?      @@      �?      @      �?      �?              �?      �?                       @              =@      @      @              �?      @      @              @      @             �E@      G@      4@       @      4@      �?      �?      �?              �?      �?              3@                      �?      7@      F@      2@      1@      @              .@      1@      �?       @      �?      @              @      �?      �?      �?                      �?              @      ,@      "@      *@      @      (@      @      @      @      �?      @               @      �?      �?              �?      �?              @              @              �?      @      �?       @      �?                       @              �?      �?      @      �?                      @      @      ;@              4@      @      @       @      @              @       @              @      @              @      @             0p@     �Q@      *@      9@      *@      @      @      @       @              �?      @      �?                      @      $@       @      $@      �?      @              @      �?      �?      �?      �?                      �?       @                      �?              2@     �n@      G@      N@      ?@      .@             �F@      ?@      @      1@      @      1@              1@      @              �?             �C@      ,@               @     �C@      (@      B@      @      7@      @      4@              @      @      @      �?      @                      �?               @      *@              @      "@      �?       @              @      �?      @              @      �?      �?              �?      �?               @      �?       @                      �?     @g@      .@     �f@      *@     �f@      $@     �e@      @     �e@      @     @R@      @      O@      �?      @      �?      @                      �?      M@              &@       @      @              @       @       @       @               @       @              @             �X@                       @      &@      @      &@       @      @       @       @       @      �?       @      �?                       @      �?              @              @                      @              @      @       @      @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJu�7hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKŅ�h��B+         F       	          ����?p�Vv���?�           ��@       3                    �?X~�pX��?�            �v@              
             �?BA�V�?�            �r@       	                    �?      �?0             R@                          �Q@      �?	             (@������������������������       �                      @                           �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@
              	          833�?R���Q�?'             N@                          `c@p���?             I@������������������������       �                    �F@                          �d@z�G�z�?             @                          �k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?z�G�z�?             $@                          q@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?       (                    �? d�=��?�            @l@                           P@�MWl��?#            �L@������������������������       �                     @                          �c@8�Z$���?             J@������������������������       �                    �B@       '                   xq@��S���?
             .@                           �?�q�q�?	             (@������������������������       �                     �?       &                    @K@�eP*L��?             &@        %                   @b@�q�q�?             "@!       "                   �e@؇���X�?             @������������������������       �                     @#       $                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @)       *                    �J@PA��ڡ?k             e@������������������������       �        C             \@+       2                   pg@�}�+r��?(            �L@,       -                   Hp@h�����?'             L@������������������������       �                    �F@.       /                    �?"pc�
�?	             &@������������������������       �                     @0       1                   Xp@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?4       E                   Pd@��y�:�?,            �P@5       >       
             �?^l��[B�?'             M@6       9                    �? >�֕�?            �A@7       8                    \@r�q��?             @������������������������       �                     �?������������������������       �                     @:       ;                    �O@XB���?             =@������������������������       �                     ;@<       =                   `a@      �?              @������������������������       �                     �?������������������������       �                     �??       @                    �?
;&����?             7@������������������������       �                     @A       B                    �?�t����?	             1@������������������������       �                     @C       D                   �h@�q�q�?             (@������������������������       �                     @������������������������       �                     @������������������������       �                     "@G       �                    �?�zц��?�            w@H       ]                    �?�B�3�?�            `p@I       V                   pp@������?            �F@J       Q                    �?���Q��?             9@K       P       	          033@X�Cc�?             ,@L       M                    �?ףp=
�?             $@������������������������       �                     @N       O       
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @R       S                    b@�C��2(�?             &@������������������������       �                      @T       U                    �J@�q�q�?             @������������������������       �                     �?������������������������       �                      @W       X                    @I@ףp=
�?             4@������������������������       �                     �?Y       \                    �?�}�+r��?             3@Z       [       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             0@^       y                    �?$Nz�{�?�             k@_       `       	          033�?xJ��b,�?k            @c@������������������������       �        "             I@a       r       
             �?ܾ�z�<�?I             Z@b       q                    �M@      �?C             X@c       f                   �Z@�j��b�?*            �M@d       e                    �?      �?             @������������������������       �                      @������������������������       �                      @g       n                    @M@,�+�C�?'            �K@h       m                    \@���J��?%            �I@i       j                    �K@؇���X�?             @������������������������       �                     @k       l       	             @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      F@o       p       
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �B@s       v                    �O@      �?              @t       u                   `l@z�G�z�?             @������������������������       �                     @������������������������       �                     �?w       x                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?z       �       	          ����?�? Da�?(            �O@{       �                   �`@      �?             4@|       �                   �X@�r����?	             .@}       �                   0a@���Q��?             @~                          (q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                   �]@���Q��?             @������������������������       �                      @������������������������       �                     @�       �       	          ����?Du9iH��?            �E@�       �                    �?�r����?             .@�       �                     O@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?$�q-�?             *@�       �       
             �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   P`@h�����?             <@�       �                   @]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     9@�       �       
             �?�"��61�?I            �Z@�       �                   �s@��qC�?6            �S@�       �                    @L@|�i���?4             S@�       �       	             @�xGZ���?            �A@�       �                    �?և���X�?             <@������������������������       �                     &@�       �                    �?�t����?             1@�       �                    �?և���X�?             @������������������������       �                     @�       �                    �K@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �_@ףp=
�?	             $@�       �                   �\@z�G�z�?             @������������������������       �                     @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �R@��r._�?            �D@�       �                   pb@�ݜ�?            �C@�       �                   P`@�FVQ&�?            �@@�       �                    `@�<ݚ�?	             "@������������������������       �                     @������������������������       �                      @������������������������       �                     8@�       �                    �?      �?             @�       �                     P@���Q��?             @������������������������       �                      @�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       	          ���@��X��?             <@�       �                    �?�㙢�c�?             7@�       �                    �?�}�+r��?             3@�       �                     M@��S�ۿ?
             .@������������������������       �                     $@�       �                   �c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �P@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK�KK��ha�BP       @t@     �y@     @o@     �\@     �l@     �Q@      2@      K@      "@      @               @      "@      �?              �?      "@              "@     �I@      �?     �H@             �F@      �?      @      �?      �?              �?      �?                      @       @       @       @      �?       @                      �?              �?     @j@      0@      F@      *@              @      F@       @     �B@              @       @      @      @      �?              @      @      @      @      @      �?      @               @      �?              �?       @                       @               @              @     �d@      @      \@              K@      @      K@       @     �F@              "@       @      @              @       @               @      @                      �?      6@     �F@      *@     �F@       @     �@@      �?      @      �?                      @      �?      <@              ;@      �?      �?      �?                      �?      &@      (@      @              @      (@              @      @      @              @      @              "@             �R@     pr@      =@      m@      (@     �@@      $@      .@      "@      @      "@      �?      @              @      �?              �?      @                      @      �?      $@               @      �?       @      �?                       @       @      2@      �?              �?      2@      �?       @               @      �?                      0@      1@      i@      "@      b@              I@      "@     �W@      @     �V@      @     �J@       @       @       @                       @      @     �I@      �?      I@      �?      @              @      �?      @      �?                      @              F@      @      �?              �?      @                     �B@      @      @      �?      @              @      �?               @      �?       @                      �?       @     �K@      @      .@       @      *@       @      @       @      �?       @                      �?               @              $@      @       @               @      @              @      D@       @      *@      �?      �?              �?      �?              �?      (@      �?      @              @      �?                      @      �?      ;@      �?       @               @      �?                      9@     �F@      O@      :@     �J@      7@     �J@      0@      3@      0@      (@      &@              @      (@      @      @      @              �?      @              @      �?              �?      "@      �?      @              @      �?      �?              �?      �?                      @              @      @      A@      @      A@       @      ?@       @      @              @       @                      8@      @      @      @       @       @              �?       @      �?                       @              �?       @              @              3@      "@      3@      @      2@      �?      ,@      �?      $@              @      �?      @                      �?      @              �?      @      �?                      @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��!XhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKՅ�h��B�.         v                    �?U�ք�?�           ��@       e                    �?n�����?           @z@       .       
             �?do@I�l�?�            �t@       +                    �?^H���+�?L            �[@                           �?�������?G            �Y@              	          ����?fP*L��?              F@������������������������       �                     ,@              	          ����?�������?             >@	       
       	          ����?r�q��?             @������������������������       �                     @                          pd@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           e@�8��8��?             8@                          �c@�nkK�?             7@������������������������       �                     �?������������������������       �                     6@������������������������       �                     �?                          �f@TV����?'            �M@                           @G@�8��8��?             (@                           _@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@                          �l@JJ����?            �G@������������������������       �                     ,@       *                   0f@�q�q�?            �@@       '                     P@¦	^_�?             ?@       $                    �?���B���?             :@                           �?�q�q�?             @������������������������       �                     @        !                   Pm@�q�q�?             @������������������������       �                     �?"       #                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?%       &                   �r@P���Q�?
             4@������������������������       �        	             3@������������������������       �                     �?(       )                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @,       -       	             �?      �?              @������������������������       �                      @������������������������       �                     @/       d                   h@      �?�             l@0       c       	             @X�*��?�            �k@1       \                   �t@��s97�?�            �k@2       W       	          ����?�V���?�            �j@3       H                   Pb@Xʃ=��?�            �i@4       A                    ]@��v$���?w            �f@5       >                   �e@@4և���?             <@6       =                    �? ��WV�?             :@7       <                    �F@�C��2(�?             &@8       9                   �[@z�G�z�?             @������������������������       �                     �?:       ;                   pb@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        	             .@?       @                   @f@      �?              @������������������������       �                     �?������������������������       �                     �?B       G                    �? u�z\A�?f            `c@C       F                    �?h�����?             <@D       E                   Pf@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     9@������������������������       �        R            �_@I       N                    @L@��s����?             5@J       M                    �D@��S�ۿ?             .@K       L                    m@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@O       V                    �Q@      �?             @P       Q                    �?���Q��?             @������������������������       �                     �?R       S                    @      �?             @������������������������       �                      @T       U       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?X       Y                   `o@"pc�
�?             &@������������������������       �                      @Z       [                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @]       ^                    �?�q�q�?             @������������������������       �                     �?_       `                   @`@���Q��?             @������������������������       �                     �?a       b                   �u@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     �?f       s       
             �?ܻ�yX7�?4            @U@g       r                   �x@����˵�?#            �M@h       q                   �`@XB���?"             M@i       p       	          ���@�>����?             ;@j       o                    @L@ ��WV�?             :@k       n                    �?@4և���?             ,@l       m                   �j@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �                     �?������������������������       �                     ?@������������������������       �                     �?t       u                   �O@�n_Y�K�?             :@������������������������       �                     $@������������������������       �        
             0@w       �                    �?JN�#:�?�            �s@x       �                   Pd@�R����?�            @n@y       �                   pf@H0sE�d�?�             l@z       �       
             �?�����?�            �k@{       �                   0a@�"P��?{            �h@|       �                   Pr@x��-�?c            �c@}       �                   p`@5�wAd�?S            �`@~       �                   @\@@4և���?)             L@       �                   �i@     ��?             0@������������������������       �                      @�       �                   �^@      �?              @������������������������       �                     @�       �                    �?      �?             @�       �                    @L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    \@�(\����?             D@�       �       	             �?ףp=
�?             $@�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     >@�       �                    �?�(�Tw�?*            �S@�       �                    l@p���?             I@������������������������       �                    �@@�       �                   �[@�IєX�?             1@�       �                   �m@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     <@�       �                   �^@z�G�z�?             9@�       �       
             �?�n_Y�K�?             *@������������������������       �                     @�       �       	             �?z�G�z�?             $@�       �                   �Y@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     (@�       �                   �m@8�Z$���?            �C@�       �                    �?�z�G��?             4@������������������������       �                     @�       �                   Pm@@�0�!��?             1@�       �                   �Z@��S�ۿ?             .@������������������������       �                     �?������������������������       �        
             ,@������������������������       �                      @������������������������       �                     3@�       �                    �?�q�q�?             8@������������������������       �                      @�       �                    �G@�GN�z�?             6@������������������������       �                      @�       �       	          ����?R���Q�?             4@�       �                    �I@�<ݚ�?             "@������������������������       �                     �?�       �                   �l@      �?              @�       �                    @O@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   `b@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     @������������������������       �                     1@�       �                    �?�q�q�?2             R@�       �       
             �?6C�z��?(            �L@�       �       	          @33�?��Sݭg�?            �C@������������������������       �                     @�       �                   �c@     ��?             @@������������������������       �                     (@�       �                   �a@      �?             4@�       �                   �l@�	j*D�?
             *@������������������������       �                     @�       �                   �r@�q�q�?             @�       �                   �b@z�G�z�?             @������������������������       �                     @�       �                    e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     �?�       �                    �?r�q��?             @������������������������       �                     @�       �                   `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     2@�       �                   �d@�r����?
             .@������������������������       �        	             *@������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK�KK��ha�BP        t@     �y@     �p@      c@      o@     �U@     �C@      R@     �@@     �Q@      @     �B@              ,@      @      7@      @      �?      @               @      �?       @                      �?       @      6@      �?      6@      �?                      6@      �?              :@     �@@      �?      &@      �?       @      �?                       @              "@      9@      6@      ,@              &@      6@      "@      6@      @      5@      @       @      @              �?       @              �?      �?      �?      �?                      �?      �?      3@              3@      �?              @      �?      @                      �?       @              @       @               @      @             @j@      ,@     @j@      *@     @j@      &@     �i@      "@     �h@      @     �f@      @      :@       @      9@      �?      $@      �?      @      �?      �?              @      �?      @                      �?      @              .@              �?      �?              �?      �?             @c@      �?      ;@      �?       @      �?              �?       @              9@             �_@              1@      @      ,@      �?      @      �?              �?      @              &@              @      @      @       @              �?      @      �?       @              �?      �?              �?      �?                      �?      "@       @       @              �?       @      �?                       @      @       @      �?              @       @      �?               @       @               @       @                       @              �?      3@     �P@      @      L@       @      L@       @      9@      �?      9@      �?      *@      �?      $@              $@      �?                      @              (@      �?                      ?@      �?              0@      $@              $@      0@              K@     @p@      8@     @k@      8@      i@      5@      i@      0@     �f@      $@     �b@      @      `@      @      J@      @      *@               @      @      @              @      @      �?      �?      �?              �?      �?               @              �?     �C@      �?      "@      �?       @               @      �?                      @              >@      �?     @S@      �?     �H@             �@@      �?      0@      �?      @      �?                      @              "@              <@      @      4@      @       @      @               @       @       @       @               @       @                      @              (@      @     �@@      @      ,@      @              @      ,@      �?      ,@      �?                      ,@       @                      3@      @      3@               @      @      1@       @              @      1@       @      @      �?              �?      @      �?      @      �?                      @              @      �?      $@              $@      �?              @                      1@      >@      E@      <@      =@      $@      =@              @      $@      6@              (@      $@      $@      "@      @      @               @      @      �?      @              @      �?      �?      �?                      �?      �?              �?      @              �?      �?      @              @      �?       @      �?                       @      2@               @      *@              *@       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJC�NhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK酔h��B�2         �                    �?4�5����?�           ��@       9                    �?����&�?           Py@       ,                    �?ZSu6��?i             d@       )       	          ����?o�����?K             ]@              
             �?և���X�??            �X@                          �c@�����?             C@              	          ����?�n`���?             ?@������������������������       �                     3@	       
       	          ����?      �?             (@������������������������       �                     @                           @Q@؇���X�?             @������������������������       �                     @������������������������       �                     �?                          0a@؇���X�?             @������������������������       �                     @                          xu@      �?              @������������������������       �                     �?������������������������       �                     �?       $       	          ����?������?'             N@                           �?:	��ʵ�?            �F@                          0j@      �?	             (@������������������������       �                     @                           @F@      �?              @������������������������       �                     �?                          �b@؇���X�?             @������������������������       �                     @������������������������       �                     �?                           @D@�FVQ&�?            �@@                          �e@      �?             @������������������������       �                     @������������������������       �                     �?        !                    b@XB���?             =@������������������������       �                     6@"       #                   �b@؇���X�?             @������������������������       �                     �?������������������������       �                     @%       &                   �^@��S���?	             .@������������������������       �                     @'       (                    �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @*       +       
             �?�X�<ݺ?             2@������������������������       �                     1@������������������������       �                     �?-       8                    @M@z�G�z�?            �F@.       5                   ``@8^s]e�?             =@/       0       	          ����?�㙢�c�?             7@������������������������       �        	             ,@1       4       	             �?X�<ݚ�?             "@2       3                    @E@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @6       7                    @I@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@:       o       
             �?�L�� ��?�            �n@;       h                    �?�M��?�            �i@<       =                   Pf@�q��/��?a            `b@������������������������       �                     9@>       ?                   �f@f>�cQ�?N            �^@������������������������       �                      @@       M                    �G@�r����?M             ^@A       H                    �F@�t����?             1@B       C                    �?�C��2(�?             &@������������������������       �                      @D       G                   �j@�����H�?             "@E       F       	              @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @I       J                    �?�q�q�?             @������������������������       �                      @K       L                    �?      �?             @������������������������       �                      @������������������������       �                      @N       [       	          ����?���z�k�?B            �Y@O       V                   �[@�c�Α�?             =@P       U                    @K@��S���?
             .@Q       T                    �I@�����H�?             "@R       S                   �Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @W       Z                   `^@@4և���?	             ,@X       Y                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @\       c                   �_@xL��N�?/            �R@]       b                    �?؇���X�?
             ,@^       a       	          `ff�?$�q-�?	             *@_       `                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?d       e                    @M@ �.�?Ƞ?%             N@������������������������       �                     F@f       g                   �b@      �?             0@������������������������       �                     .@������������������������       �                     �?i       j                   �r@ _�@�Y�?&             M@������������������������       �        "             J@k       l       	             �?r�q��?             @������������������������       �                     @m       n       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?p                          @b@�(�Tw��?            �C@q       z                   �d@؇���X�?             <@r       y                    �?HP�s��?             9@s       x       	          033�?�r����?             .@t       u                   �o@@4և���?
             ,@������������������������       �                      @v       w                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@{       |                    a@�q�q�?             @������������������������       �                     �?}       ~                   pf@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �\@���|���?             &@������������������������       �                     @������������������������       �                     @�       �                    �?������?�            �t@�       �                    �?f��N�&�?�            �q@�       �                    @L@�ۓ����?�            `n@�       �                   d@(S��C��?{             h@�       �                    �?      �?             ,@������������������������       �                     @�       �       	          ����?�z�G��?             $@�       �                    �?���Q��?             @������������������������       �                      @�       �       	          ������q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       
             �?���oY��?o            `f@�       �                     J@h+�v:�?             A@�       �                    �?r�q��?             8@�       �                   `b@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �       
             �?������?	             .@������������������������       �                      @�       �                   �k@�	j*D�?             *@������������������������       �                     @�       �       	          ����?ףp=
�?             $@������������������������       �                     @�       �                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                   �g@@��t��?]             b@�       �                    @G@@Tn�kq�?\            �a@������������������������       �        0            �T@�       �                   n@ �.�?Ƞ?,             N@������������������������       �                     @@�       �                    �G@h�����?             <@�       �                   �]@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@������������������������       �                      @�       �                   �u@��H�}�?#             I@�       �                    �?֭��F?�?!            �G@�       �                   ``@�t����?             1@�       �                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `_@��S�ۿ?
             .@�       �       	          ����?�q�q�?             @�       �                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                   �c@��S���?             >@�       �       	          ����?���|���?             6@�       �                    `@��S�ۿ?             .@�       �                   �m@      �?             @�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        	             &@������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   �_@�G�z��?             D@�       �                   P`@�C��2(�?             6@�       �       
             �?z�G�z�?             $@�       �                   �_@�����H�?             "@������������������������       �                     @�       �                    s@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                   �f@�����H�?             2@�       �                    �J@�IєX�?             1@������������������������       �                     (@�       �                    �K@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �       	            �?nM`����?             G@�       �       	          ���ٿz�G�z�?             .@������������������������       �                     �?�       �       	          ����?؇���X�?             ,@�       �                   �W@z�G�z�?             $@������������������������       �                     �?�       �                    �?�����H�?             "@������������������������       �                     @�       �       
             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �b@�חF�P�?             ?@������������������������       �                     6@�       �       
             �?X�<ݚ�?             "@������������������������       �                      @�       �                    �?և���X�?             @�       �                    e@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�t�b�m     h�h*h-K ��h/��R�(KK�KK��ha�B�       �t@     y@      X@     Ps@     �P@     �W@     �L@     �M@      L@      E@      (@      :@      @      9@              3@      @      @      @              �?      @              @      �?              @      �?      @              �?      �?              �?      �?              F@      0@     �B@       @      @      @              @      @       @              �?      @      �?      @                      �?      ?@       @      @      �?      @                      �?      <@      �?      6@              @      �?              �?      @              @       @              @      @       @               @      @              �?      1@              1@      �?              "@      B@      "@      4@      @      3@              ,@      @      @      @      �?              �?      @                      @      @      �?              �?      @                      0@      >@     �j@      3@     @g@      2@      `@              9@      2@      Z@       @              0@      Z@      @      (@      �?      $@               @      �?       @      �?       @               @      �?                      @      @       @       @               @       @               @       @              &@      W@       @      5@      @       @      �?       @      �?       @               @      �?                      @      @              �?      *@      �?      @              @      �?                       @      @     �Q@       @      (@      �?      (@      �?      �?              �?      �?                      &@      �?              �?     �M@              F@      �?      .@              .@      �?              �?     �L@              J@      �?      @              @      �?      �?      �?                      �?      &@      <@      @      8@       @      7@       @      *@      �?      *@               @      �?      @              @      �?              �?                      $@       @      �?      �?              �?      �?              �?      �?              @      @              @      @             �m@      W@     �k@     �O@     @i@     �D@     @e@      7@      @      @      @              @      @      @       @       @              �?       @      �?                       @              @     `d@      0@      5@      *@      &@      *@      @       @      @                       @      @      &@               @      @      "@      @              �?      "@              @      �?       @      �?                       @      $@             �a@      @     �a@      �?     �T@             �M@      �?      @@              ;@      �?      @      �?              �?      @              6@                       @      @@      2@      =@      2@      .@       @      �?      �?              �?      �?              ,@      �?       @      �?      �?      �?      �?                      �?      �?              (@              ,@      0@      ,@       @      ,@      �?      @      �?      �?      �?      �?                      �?       @              &@                      @               @      @              2@      6@       @      4@       @       @      �?       @              @      �?      @              @      �?              �?                      (@      0@       @      0@      �?      (@              @      �?              �?      @                      �?      1@      =@      (@      @              �?      (@       @       @       @              �?       @      �?      @              @      �?              �?      @              @              @      :@              6@      @      @       @              @      @       @      @       @                      @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�R�[hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK兔h��B2         d       	          ����?6������?�           ��@              
             �?��_���?�             w@                          ph@�4�M�f�?@            �Y@������������������������       �                     D@              	          ����?V��z4�?%             O@                          �c@X�EQ]N�?            �E@                          �`@      �?             @@������������������������       �        
             ,@	                           �?�X�<ݺ?	             2@
                          0a@$�q-�?             *@                          �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     @                          `]@���|���?             &@������������������������       �                     @                          0e@z�G�z�?             @������������������������       �                     @                          �l@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?�d�����?             3@                          �d@�q�q�?	             (@              	          833�?      �?              @������������������������       �                      @              
             �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @        !       	             �(��R%��?�            �p@������������������������       �                      @"       G                    �?��U�=��?�            �p@#       ,                   @E@��H�}�?0            �R@$       %                    �?8�Z$���?	             *@������������������������       �                     @&       +       	          @33�?����X�?             @'       *                    �?���Q��?             @(       )                   �]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @-       :                    �?r֛w���?'             O@.       9                   �^@�t����?             1@/       8                   `\@      �?             $@0       7                    q@      �?              @1       6                   �c@���Q��?             @2       5       	          @33�?�q�q�?             @3       4                    �H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @;       D                   �b@�:�^���?            �F@<       =                   �c@������?            �D@������������������������       �                     @@>       C                   Pd@�<ݚ�?             "@?       B                    �?�q�q�?             @@       A                    `@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @E       F                   �d@      �?             @������������������������       �                      @������������������������       �                      @H       K                   `Q@ 7���B�?z            �g@I       J                    �?�z�G��?             $@������������������������       �                     @������������������������       �                     @L       S                    @L@P�p�_�?u            `f@M       R                    �G@@�`%���?^            `b@N       O                    @G@ �й���?0            @R@������������������������       �        .            �Q@P       Q                    o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        .            �R@T       W                    �L@     ��?             @@U       V                    �?      �?              @������������������������       �                     �?������������������������       �                     �?X       a                    @��S�ۿ?             >@Y       Z                    �? ��WV�?             :@������������������������       �        	             *@[       \                   Pc@$�q-�?	             *@������������������������       �                     @]       ^                   ht@r�q��?             @������������������������       �                     @_       `                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?b       c                    �?      �?             @������������������������       �                     �?������������������������       �                     @e       �       
             �?xƅd�?�            �v@f       �                   pb@�=�y.�?�            �s@g       �       	          `ff�?��a��?�            �n@h       y                    �?�z����?W            @`@i       n                   `\@�q�q�?             B@j       k                   ``@      �?
             0@������������������������       �                     @l       m                   �t@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @o       x                    �?      �?             4@p       q                    _@����X�?             ,@������������������������       �                     @r       s                   �[@և���X�?             @������������������������       �                      @t       w       	             �?���Q��?             @u       v       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @z       �                    @�*/�8V�?>            �W@{       �                   @e@��a�n`�?=            @W@|       �                   `_@������?:            @V@}       �       	          ����?(;L]n�?&             N@~                          �Z@HP�s��?             9@������������������������       �                     "@�       �                    �?      �?             0@�       �                    \@@4և���?	             ,@������������������������       �                     �?������������������������       �                     *@�       �                   `b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �A@�       �                    �?д>��C�?             =@������������������������       �                     @�       �       	          ����?��<b���?             7@�       �                    �?�q�q�?             "@������������������������       �                     �?�       �                   �\@      �?              @������������������������       �                     �?�       �       	          033�?؇���X�?             @������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                     L@؇���X�?
             ,@������������������������       �                     $@�       �                    `@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?�       �                   @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �U@io8�?C             ]@������������������������       �                     �?�       �                   �[@P���Q�?B            �\@������������������������       �                    �C@�       �                    �?�˹�m��?0             S@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @�       �                    _@hA� �?*            �Q@�       �                   �\@@�0�!��?	             1@������������������������       �                     @������������������������       �                     ,@������������������������       �        !            �J@�       �                    �?T�iA�?$            �Q@�       �                    �?JJ����?            �G@�       �       	          `ff @����X�?             ,@������������������������       �                     $@������������������������       �                     @�       �                    �?���|���?            �@@�       �                    @L@d}h���?             ,@�       �                   �e@և���X�?             @�       �                   Pl@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	          ����?�\��N��?
             3@������������������������       �                     @�       �                   �f@����X�?             ,@�       �                    �E@�θ�?             *@������������������������       �                     �?�       �                   pd@r�q��?             (@�       �                   �g@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   �f@8����?             7@�       �       	          033�?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �Z@���y4F�?             3@�       �                   �Y@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    q@      �?	             0@������������������������       �                     (@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    ]@� �	��?$             I@������������������������       �                     @�       �                    �?F�����?             �F@�       �                    �?d}h���?             <@������������������������       �                     "@�       �                    d@�����?             3@�       �                   `U@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                   �l@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?ҳ�wY;�?             1@�       �                    �?      �?
             (@�       �                   @`@      �?              @������������������������       �                     �?�       �                    S@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK�KK��ha�BP       �t@     �x@      o@     �]@      3@     �T@              D@      3@     �E@      @      C@      �?      ?@              ,@      �?      1@      �?      (@      �?      @      �?                      @              "@              @      @      @              @      @      �?      @              �?      �?      �?                      �?      ,@      @      @      @      @      @       @              �?      @      �?                      @      @              @             �l@      B@               @     �l@      A@      H@      ;@       @      &@              @       @      @       @      @       @       @       @                       @              �?               @      G@      0@      @      (@      @      @      @      @      @       @      �?       @      �?      �?              �?      �?                      �?       @                      @       @                      @     �D@      @     �C@       @      @@              @       @      �?       @      �?      �?      �?                      �?              �?      @               @       @               @       @             �f@      @      @      @              @      @             �e@      @     @b@      �?      R@      �?     �Q@              �?      �?              �?      �?             �R@              =@      @      �?      �?              �?      �?              <@       @      9@      �?      *@              (@      �?      @              @      �?      @              �?      �?      �?                      �?      @      �?              �?      @             �U@     �q@      M@      p@      =@      k@      6@      [@      (@      8@       @      ,@              @       @      @              @       @              $@      $@      $@      @      @              @      @               @      @       @      �?       @      �?                       @       @                      @      $@      U@      "@      U@      @     �T@       @      M@       @      7@              "@       @      ,@      �?      *@      �?                      *@      �?      �?              �?      �?                     �A@      @      8@              @      @      2@      @      @      �?               @      @      �?              �?      @               @      �?      @              @      �?               @      (@              $@       @       @       @                       @       @       @              �?       @      �?              �?       @              �?              @     @[@      �?              @     @[@             �C@      @     �Q@      @      @              @      @              @     �P@      @      ,@      @                      ,@             �J@      =@     �D@      6@      9@      $@      @      $@                      @      (@      5@      @      &@      @      @      �?      @      �?                      @       @                      @      "@      $@      @              @      $@      @      $@      �?               @      $@       @      @              @       @                      @      �?              @      0@      @      �?              �?      @              @      .@       @      �?              �?       @               @      ,@              (@       @       @               @       @              <@      6@              @      <@      1@      6@      @      "@              *@      @      "@      �?              �?      "@              @      @              @      @              @      &@      @      @       @      @      �?              �?      @      �?                      @      @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�v}hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B�(         r                    �?U�ք�?�           ��@                           �?~e�.y�?
            z@                          �Q@d�.����?K            @^@������������������������       �                     @              
             �?t��%�?H            �\@                           �?��R[s�?            �A@                          `X@     ��?             @@������������������������       �                      @	                           �?�r����?             >@
                          �a@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     7@������������������������       �                     @                          @c@�(\����?4             T@������������������������       �        0             R@                           �?      �?              @������������������������       �                      @������������������������       �                     @       #                   �_@�?ȇ�p�?�            pr@                           �?j�'�=z�?)            �P@              
             �?�e����?            �C@              	          `ff�?�>4և��?             <@������������������������       �                     (@                          `_@     ��?	             0@������������������������       �                     @                          @`@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �        
             &@               
             �? 7���B�?             ;@������������������������       �        
             0@!       "                    @I@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@$       g                    @P�����?�            �l@%       ^       	          `ff�?��H.�!�?�             i@&       +                    P@�&�5y�?}            @g@'       *       	          �����@4և���?             ,@(       )       	          ���ٿ      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             (@,       M                   xp@p����?q            �e@-       F       	          ����?     ��?T             `@.       5                   �[@X�
����?K             ]@/       0                    �?      �?             8@������������������������       �                     @1       4                   0n@����X�?
             5@2       3       
             �?�t����?             1@������������������������       �                      @������������������������       �                     .@������������������������       �                     @6       A       	            �?���.�6�??             W@7       <       
             �?��`qM|�?8            �T@8       ;                    �?և���X�?             @9       :                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @=       >                   �b@�"w����?4             S@������������������������       �        1            @Q@?       @                   �c@؇���X�?             @������������������������       �                     �?������������������������       �                     @B       C                   @l@�<ݚ�?             "@������������������������       �                     @D       E                     M@�q�q�?             @������������������������       �                      @������������������������       �                     �?G       J                    �J@�q�q�?	             (@H       I                   �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?K       L                   @^@؇���X�?             @������������������������       �                     �?������������������������       �                     @N       S                   �p@8�A�0��?             F@O       P                   �c@؇���X�?             @������������������������       �                     @Q       R                    �?      �?              @������������������������       �                     �?������������������������       �                     �?T       Y                    �?4�B��?            �B@U       X                    s@���!pc�?             &@V       W                   `q@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @Z       [                   �`@8�Z$���?             :@������������������������       �                      @\       ]                    \@�8��8��?             8@������������������������       �                      @������������������������       �                     6@_       d                    `@����X�?
             ,@`       a                   �l@"pc�
�?             &@������������������������       �                      @b       c                   �o@�q�q�?             @������������������������       �                      @������������������������       �                     �?e       f                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @h       q       
             �?����"�?             =@i       p                    �P@"pc�
�?             6@j       o                    �?ףp=
�?             4@k       n                   �m@����X�?             @l       m                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@������������������������       �                      @������������������������       �                     @s       t                   �U@��Dl<�?�            �s@������������������������       �                     @u       �       
             �?����X��?�            �s@v       �                    @G@TY��&\�?�            �p@w       x                    �?�GN�z�?             F@������������������������       �                     @y       �                    �?��r._�?            �D@z       {                   �h@z�G�z�?            �A@������������������������       �                     0@|       }                   �`@p�ݯ��?             3@������������������������       �                     @~                           �A@�q�q�?             (@������������������������       �                      @�       �                    �E@�z�G��?             $@������������������������       �                     @�       �       	             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    a@�2�~w�?�            �k@�       �                    Z@�����?g            `e@������������������������       �                     F@�       �                   P`@�m(']�?O            �_@�       �                    �?������?            �B@�       �                   @s@r�q��?             8@�       �                   �d@�C��2(�?             6@������������������������       �                     *@�       �                   �Z@�<ݚ�?             "@������������������������       �                     �?�       �       	             �?      �?              @�       �                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �        
             *@�       �                    �R@�E�����?4            �V@������������������������       �        3            @V@������������������������       �                     �?�       �                   0a@ZՏ�m|�?!            �H@������������������������       �                      @�       �       	          ����?��E�B��?             �G@������������������������       �        
             ,@�       �                    �?"pc�
�?            �@@�       �                    @K@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �j@�>����?             ;@�       �                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     4@�       �                   �]@Np�����?             �I@������������������������       �                     "@�       �                    �?�D����?             E@�       �                   Pd@�f7�z�?             =@�       �                     M@`�Q��?             9@�       �                   �_@ףp=
�?             $@�       �                   @a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	          033�?��S���?	             .@�       �                   �c@���!pc�?             &@�       �                    �?և���X�?             @������������������������       �                      @�       �                     N@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     *@�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�        t@     �y@     �p@      b@      Z@      1@              @      Z@      &@      :@      "@      :@      @               @      :@      @      @      @      @                      @      7@                      @     �S@       @      R@              @       @               @      @             �d@      `@      1@     �H@      0@      7@      @      7@              (@      @      &@              @      @      @      @                      @      &@              �?      :@              0@      �?      $@      �?                      $@     �b@     �S@     `a@     �N@     �`@     �I@      �?      *@      �?      �?              �?      �?                      (@     �`@      C@      [@      4@     @Y@      .@      .@      "@              @      .@      @      .@       @               @      .@                      @     �U@      @     �S@      @      @      @      @      �?              �?      @                       @     �R@      �?     @Q@              @      �?              �?      @              @       @      @              �?       @               @      �?              @      @      �?      @              @      �?              @      �?              �?      @              :@      2@      �?      @              @      �?      �?      �?                      �?      9@      (@      @       @      �?       @      �?                       @       @              6@      @               @      6@       @               @      6@              @      $@       @      "@               @       @      �?       @                      �?       @      �?              �?       @              &@      2@      @      2@       @      2@       @      @       @      �?              �?       @                      @              *@       @              @             �I@     �p@      @              H@     �p@      7@      n@      $@      A@      @              @      A@      @      <@              0@      @      (@              @      @      @               @      @      @      @               @      @              @       @                      @      *@     �i@      @     �d@              F@      @     �^@      @     �@@      @      4@       @      4@              *@       @      @      �?              �?      @      �?       @      �?                       @              @       @                      *@      �?     @V@             @V@      �?               @     �D@       @              @     �D@              ,@      @      ;@      @       @      @                       @       @      9@       @      @              @       @                      4@      9@      :@              "@      9@      1@      (@      1@       @      1@      �?      "@      �?       @               @      �?                      @      @       @      @       @      @      @       @              �?      @      �?                      @              @      @              @              *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJg}�XhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B�5         �                    �?0����?�           ��@       A       
             �?�ua��?           @{@              	          ����?n2�`���?b            `c@                           �?�C��2(�?            �K@������������������������       �                     D@       	                    @E@�q�q�?             .@                           �?      �?             @������������������������       �                     @������������������������       �                     �?
                           �?"pc�
�?	             &@������������������������       �                     �?                          �c@ףp=
�?             $@������������������������       �                     @                          �`@      �?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           �?Fx$(�?D             Y@                           �?      �?             4@������������������������       �                     @                          `X@      �?             0@������������������������       �                     �?������������������������       �                     .@       @                   �t@���Q8�?5             T@       5                   �`@      �?3             S@       *                   Pl@8�$�>�?            �E@       #                   �^@      �?             8@                           �?z�G�z�?             $@������������������������       �                     @                           �a@���Q��?             @������������������������       �                      @!       "                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?$       %       	             �?����X�?	             ,@������������������������       �                      @&       '                    _@�q�q�?             @������������������������       �                     �?(       )                     O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?+       .                    �D@�S����?             3@,       -       	              @      �?              @������������������������       �                     �?������������������������       �                     �?/       4                     P@�t����?             1@0       1                    �?8�Z$���?	             *@������������������������       �                     �?2       3                    `@r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     @6       ?                    �?<���D�?            �@@7       <                    @O@�<ݚ�?             2@8       ;                   0a@@4և���?
             ,@9       :                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@=       >                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             .@������������������������       �                     @B       e                    �?��L��?�            �q@C       d                    �?��It��?1            �S@D       Y                   �_@�� =[�?+             Q@E       V       	          ����?���"͏�?            �B@F       M                    �?�חF�P�?             ?@G       H                   �c@      �?              @������������������������       �                     @I       J                   �d@z�G�z�?             @������������������������       �                      @K       L                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?N       O                    �?�nkK�?             7@������������������������       �                     @P       Q                    ]@      �?             0@������������������������       �                     @R       S       	          @33�?ףp=
�?             $@������������������������       �                      @T       U       	          pff�?      �?              @������������������������       �                     �?������������������������       �                     �?W       X       	             �?�q�q�?             @������������������������       �                     @������������������������       �                      @Z       _                    �?`Jj��?             ?@[       \                   �b@      �?              @������������������������       �                     @]       ^                    �?      �?             @������������������������       �                     �?������������������������       �                     @`       a                   �b@�nkK�?             7@������������������������       �                     5@b       c                    �E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@f       �                    @��5�uԾ?�            @i@g       l                   @[@p�qG�?}             h@h       i                    �?�<ݚ�?             "@������������������������       �                     @j       k                    i@�q�q�?             @������������������������       �                     �?������������������������       �                      @m       �                     R@ ��^og�?v            �f@n       u                   �P@ k��ͫ?s            `f@o       r                    �?����X�?             @p       q                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?s       t                    �?      �?              @������������������������       �                     �?������������������������       �                     �?v                          �t@��$����?m            �e@w       ~       	          ���@ ��N8�?j             e@x       y                    @L@�E��La�?i            �d@������������������������       �        X            `a@z       }                   �_@h�����?             <@{       |                   �^@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     4@������������������������       �                     �?�       �                   @`@      �?             @������������������������       �                      @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    `R@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @M@�z�G��?             $@������������������������       �                     @�       �                    @N@���Q��?             @������������������������       �                      @�       �                     P@�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �b@�q�� �?�            �r@�       �       
             �?�A����?�            @q@�       �                    �?�cX1!��?�             o@�       �                   �s@x���cB�?v            @g@�       �                    �?t�G����?n            �e@�       �                    �?     x�?S             `@�       �                   �l@      �?             0@�       �                    �H@      �?             @������������������������       �                     �?�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@�       �                   �l@���>4ֵ?H             \@�       �                   �Z@�U�:��?'            �M@������������������������       �                      @�       �                   �[@�}�+r��?&            �L@�       �                   @[@؇���X�?             ,@������������������������       �                     "@�       �                    �J@���Q��?             @������������������������       �                     �?�       �                   �k@      �?             @������������������������       �                      @������������������������       �                      @�       �                   `_@ qP��B�?            �E@������������������������       �                     7@�       �       	          ����?P���Q�?             4@�       �       	             �?؇���X�?             @������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �        !            �J@�       �                    �?��2(&�?             F@�       �                    �?      �?             @�       �                     M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �`@ףp=
�?             D@�       �                   �X@�IєX�?             A@�       �       	             @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �_@      �?             @@������������������������       �                     �?������������������������       �                     ?@�       �                    �I@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    t@����X�?             ,@������������������������       �                     @�       �                   �t@�C��2(�?             &@�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �R@���N8�?'            �O@�       �                   �`@�g�y��?&             O@������������������������       �                     H@�       �                   0a@؇���X�?	             ,@������������������������       �                      @������������������������       �                     (@������������������������       �                     �?�       �                    �?|��?���?             ;@�       �       	          ����?r�q��?             8@�       �                   �_@�	j*D�?             *@������������������������       �                     �?�       �       	             �?      �?             (@�       �                    �?���Q��?             @������������������������       �                      @�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �b@���|���?             &@�       �                    @N@և���X�?             @�       �       	             @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �I@�q�q�?             @������������������������       �                     �?�       �                    @M@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @O@���|���?             6@�       �                   �^@�z�G��?             4@������������������������       �                     @�       �                    `@և���X�?
             ,@������������������������       �                      @�       �                   �j@�q�q�?             (@�       �       	             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK�KK��ha�BP        u@     �x@     r@     `b@     �E@      \@      @      I@              D@      @      $@      @      �?      @                      �?       @      "@      �?              �?      "@              @      �?      @      �?      �?      �?                      �?               @      C@      O@      .@      @              @      .@      �?              �?      .@              7@     �L@      3@     �L@      .@      <@      (@      (@       @       @              @       @      @               @       @      �?       @                      �?      $@      @       @               @      @      �?              �?      @              @      �?              @      0@      �?      �?      �?                      �?       @      .@       @      &@              �?       @      $@              $@       @                      @      @      =@      @      ,@      �?      *@      �?      @      �?                      @              $@      @      �?              �?      @                      .@      @             �n@     �A@     �L@      6@     �L@      &@      <@      "@      :@      @      @      @              @      @      �?       @               @      �?       @                      �?      6@      �?      @              .@      �?      @              "@      �?       @              �?      �?              �?      �?               @      @              @       @              =@       @      @      �?      @              @      �?              �?      @              6@      �?      5@              �?      �?              �?      �?                      &@     �g@      *@     �f@      $@      @       @      @              �?       @      �?                       @     �e@       @     �e@      @      @       @      @      �?      @                      �?      �?      �?      �?                      �?      e@      @     �d@       @     �d@      �?     `a@              ;@      �?      @      �?      @                      �?      4@                      �?      @      �?       @              �?      �?              �?      �?              �?      @              �?      �?       @               @      �?              @      @      @               @      @               @       @      �?      �?              �?      �?      �?                      �?     �G@     `o@     �@@     `n@      4@     �l@      1@      e@      *@     �c@      @     @^@       @      ,@       @       @              �?       @      �?              �?       @                      (@      @     �Z@      @      K@       @              @      K@       @      (@              "@       @      @              �?       @       @               @       @              �?      E@              7@      �?      3@      �?      @              @      �?      �?      �?                      �?              *@             �J@      @      C@       @       @       @      �?              �?       @                      �?      @      B@       @      @@      �?      �?      �?                      �?      �?      ?@      �?                      ?@       @      @       @                      @      @      $@      @              �?      $@      �?       @               @      �?                       @      @      N@       @      N@              H@       @      (@       @                      (@      �?              *@      ,@      &@      *@      @      "@      �?              @      "@      @       @       @              �?       @               @      �?                      @      @      @      @      @      @      �?      @                      �?              @      @               @      �?      �?              �?      �?              �?      �?              ,@       @      ,@      @      @               @      @               @       @      @      �?      @      �?                      @      @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ	�tlhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK˅�h��Bh,         b                    �?�+	G�?�           ��@       =       
             �?��4:���?�            Px@       <                   �e@�č����?�            �r@                          �k@�Tޫvɼ?�            �r@                           �?p�`Bh�?a            �b@              
             �?      �?	             0@������������������������       �                      @       	                   �R@؇���X�?             ,@������������������������       �                      @
                           �?�q�q�?             @������������������������       �                      @������������������������       �                     @                           �?`��(�?X            �`@������������������������       �        C            �X@                           �?@-�_ .�?            �B@              
             �?�KM�]�?	             3@                          �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@������������������������       �                     2@                          �m@���Lͩ�?b            �b@                           �G@      �?             <@������������������������       �                     @                          �_@      �?             8@������������������������       �                     1@                           �?և���X�?             @              	             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @        ;                    �R@ @|���?Q            �^@!       "                   �Q@����&!�?P            @^@������������������������       �                     �?#       2                    c@ �q�q�?O             ^@$       +       	          033@�O4R���?F            �Z@%       &                    @N@��f�{��?8            �U@������������������������       �        +            �P@'       *                    �?P���Q�?             4@(       )                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     1@,       1                    �J@P���Q�?             4@-       0                   pq@      �?             @.       /       	             @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     0@3       8       	          `ff�?d}h���?	             ,@4       5                    �N@�����H�?             "@������������������������       �                     @6       7                    �?      �?             @������������������������       �                     �?������������������������       �                     @9       :       	          `ff@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                      @>       M                   @E@�a7���?4            �U@?       @                    �G@��}*_��?             ;@������������������������       �                     @A       B                   �X@      �?             4@������������������������       �                      @C       D                    �?X�<ݚ�?
             2@������������������������       �                     �?E       L                   �a@j���� �?	             1@F       G                    [@�q�q�?             (@������������������������       �                     @H       K                    �?�<ݚ�?             "@I       J                     P@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @N       [                    �?��mo*�?$            �M@O       Z                    �?���Q��?             .@P       Q                   �b@�q�q�?             "@������������������������       �                     @R       Y       	          @33�?      �?             @S       T                    ]@���Q��?             @������������������������       �                     �?U       V                   d@      �?             @������������������������       �                      @W       X                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @\       ]                   �c@�Ra����?             F@������������������������       �                     6@^       _                   �`@�GN�z�?             6@������������������������       �                     (@`       a                   �l@      �?             $@������������������������       �                     @������������������������       �                     @c       �       	          pff�?bPD΂_�?�            �u@d       w                   �\@     |�?�             p@e       j                   �j@�G��l��?             5@f       i                    �?      �?              @g       h                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @k       t                   �`@�	j*D�?	             *@l       m                    W@z�G�z�?             $@������������������������       �                     @n       s       
             �?����X�?             @o       r                    �?      �?             @p       q                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @u       v                   @X@�q�q�?             @������������������������       �                      @������������������������       �                     �?x       �                   @g@�7��d��?�            `m@y       �       
             �?�8h
Q��?�             m@z       �                   �`@�LQ�1	�?              G@{       ~                   �a@؇���X�?             <@|       }       	          `ff�?      �?             @������������������������       �                     @������������������������       �                     @       �                    ]@���7�?             6@�       �                    �?�q�q�?             @������������������������       �                     �?�       �       	          @33�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             3@�       �                   �c@�q�q�?             2@�       �                     R@d}h���?             ,@�       �                   @a@8�Z$���?
             *@�       �                   0e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?@>ZAɥ�?q            `g@������������������������       �        #             M@�       �                    @L@���f�?N             `@�       �                   0n@@䯦s#�?@            �Z@������������������������       �        (            �M@�       �                   �n@`Ql�R�?            �G@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                    �E@�       �                    �?�㙢�c�?             7@�       �                   �p@������?	             .@�       �       	            �?      �?              @������������������������       �                      @�       �                    a@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    �?�VM�?6            @V@�       �                    �L@V{q֛w�?&             O@�       �                    �?�	j*D�?             :@������������������������       �                     *@�       �                    �?�n_Y�K�?
             *@������������������������       �                     @�       �                    �K@z�G�z�?	             $@�       �                   �\@�����H�?             "@������������������������       �                     @�       �                    @E@r�q��?             @�       �       	             @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �n@      �?             B@�       �                   Pd@��H�}�?             9@�       �                    �?�\��N��?             3@������������������������       �                      @�       �       	              @j���� �?             1@�       �                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �                   `a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                   @^@�>����?             ;@������������������������       �                     �?�       �                    �I@ ��WV�?             :@�       �       	          033�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       `t@     �y@     �R@     �s@      4@     �q@      2@     �q@      @     `b@       @      ,@               @       @      (@               @       @      @       @                      @       @     �`@             �X@       @     �A@       @      1@       @      �?       @                      �?              0@              2@      ,@      a@      @      5@      @              @      5@              1@      @      @      @       @      @                       @               @      @     �\@      @     �\@      �?              @     �\@       @      Z@      �?     @U@             �P@      �?      3@      �?       @               @      �?                      1@      �?      3@      �?      @      �?      �?      �?                      �?               @              0@      @      &@      �?       @              @      �?      @      �?                      @       @      @       @                      @      �?               @             �K@      ?@      $@      1@              @      $@      $@               @      $@       @              �?      $@      @      @      @      @               @      @       @       @       @                       @              @      @             �F@      ,@      @      "@      @      @      @              @      @      @       @              �?      @      �?       @              �?      �?      �?                      �?              �?              @     �C@      @      6@              1@      @      (@              @      @              @      @             `o@     �W@     �k@      A@      $@      &@      �?      @      �?      �?              �?      �?                      @      "@      @       @       @      @              @       @       @       @       @      �?       @                      �?              �?      @              �?       @               @      �?             �j@      7@     �j@      5@      >@      0@      8@      @      @      @              @      @              5@      �?       @      �?      �?              �?      �?              �?      �?              3@              @      (@      @      &@       @      &@      �?      �?      �?                      �?      �?      $@      �?                      $@      �?              @      �?      @                      �?     �f@      @      M@              _@      @     @Z@      �?     �M@              G@      �?      @      �?      @                      �?     �E@              3@      @      &@      @      @      @       @               @      @              @       @              @               @                       @      =@      N@      ;@     �A@      2@       @      *@              @       @      @               @       @      �?       @              @      �?      @      �?      �?      �?                      �?              @      �?              "@      ;@      "@      0@      "@      $@       @              @      $@      @      @      @                      @      �?      @              @      �?      �?              �?      �?                      @              &@       @      9@      �?              �?      9@      �?      @      �?                      @              6@�t�bub�0     hhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�ޡhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKǅ�h��B�+         x                    �?6������?�           ��@       [       	          ����?�C�"��?"           �{@                          `_@n(��"�?�            v@                           �?��
ц��?.            @P@������������������������       �        
             1@                           @K@      �?$             H@       
       
             �?r�q��?             8@       	       
             �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@              	             �?$�q-�?             *@������������������������       �        
             (@������������������������       �                     �?              
             �?�q�q�?             8@                          8w@�X�<ݺ?             2@������������������������       �                     1@������������������������       �                     �?                           @M@�q�q�?             @������������������������       �                      @                           �N@      �?             @������������������������       �                      @������������������������       �                      @       $                    �?F��ӭ��?�             r@       !                    �?�}#���?6            �T@                            �?p�|�i�?0             S@                          �r@      �?             (@                           ^@ףp=
�?             $@              
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �        )             P@"       #       
             �?և���X�?             @������������������������       �                     @������������������������       �                     @%       8       
             �?B�黀;�?�            �i@&       -       	          ����?ҳ�wY;�?            �I@'       ,                    �?��S�ۿ?             >@(       )                    �?�����?             5@������������������������       �                     &@*       +                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     "@.       7                    @O@���N8�?             5@/       0                    �G@X�Cc�?
             ,@������������������������       �                     @1       6       	          ����?X�<ݚ�?             "@2       3                    �?�q�q�?             @������������������������       �                     @4       5                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @9       D                    �?T����?c            @c@:       ;                   �b@J�8���?             =@������������������������       �                     @<       =                   `\@\X��t�?             7@������������������������       �                     @>       C                   �d@������?             1@?       B                    �?@4և���?             ,@@       A                   @f@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                     @E       V       	          pff�?0{�v��?N            @_@F       S                   xt@�7��?H            @]@G       N                   �b@�?�|�?F            �[@H       I                   Hp@�ջ����?B             Z@������������������������       �        4             S@J       K                     L@h�����?             <@������������������������       �                     :@L       M                    q@      �?              @������������������������       �                     �?������������������������       �                     �?O       R       	          @33�?����X�?             @P       Q                   @f@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?T       U                    �?      �?             @������������������������       �                     @������������������������       �                     @W       X                   �^@      �?              @������������������������       �                     @Y       Z                   �b@���Q��?             @������������������������       �                      @������������������������       �                     @\       s       	          ��� @���?>            @V@]       f                   �b@����e��?.            �P@^       e                    �?� ��1�?            �D@_       `                   pe@�	j*D�?             :@������������������������       �                     @a       b                   �a@؇���X�?             5@������������������������       �                     0@c       d                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        
             .@g       n                   �p@ �o_��?             9@h       m                   �_@@4և���?             ,@i       l       	             �?z�G�z�?             @j       k                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@o       p                    �?�eP*L��?             &@������������������������       �                     @q       r                    @I@؇���X�?             @������������������������       �                     �?������������������������       �                     @t       u                    @�nkK�?             7@������������������������       �                     4@v       w                   0`@�q�q�?             @������������������������       �                     �?������������������������       �                      @y       �       
             �?v���a�?�            @r@z       �                    �?$%j����?�            �o@{       �                    l@(L���?o            �e@|       }                   �U@ ��Ou��?3            �S@������������������������       �                      @~                          0a@p�|�i�?2             S@������������������������       �        *            �P@�       �                    �J@�z�G��?             $@�       �                    �H@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   pl@ظ�*���?<            �W@������������������������       �                     @�       �                   �l@4\�����?;            @V@�       �                    �?���Q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �a@؇���X�?7             U@�       �       	          ����?�rF���?%            �K@�       �                    �?��H�}�?             9@�       �                   @b@�E��ӭ�?             2@�       �                    �?������?             1@������������������������       �                      @�       �                    �?�r����?
             .@������������������������       �                      @�       �                   �p@8�Z$���?             *@�       �       	          433�?���Q��?             @������������������������       �                     �?�       �                   �\@      �?             @������������������������       �                     �?�       �                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    �?և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   Pa@ףp=
�?             >@�       �       	          033@ ��WV�?             :@������������������������       �                     3@�       �                   �\@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    �M@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     =@�       �                   @s@ �)���?6            @T@������������������������       �        0             R@�       �       
             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �       	          ����?Hث3���?            �C@�       �                   @`@�<ݚ�?             2@�       �                    �I@      �?             @������������������������       �                      @������������������������       �                      @�       �                   d@؇���X�?             ,@������������������������       �                      @�       �                    h@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �D@���N8�?             5@������������������������       �                      @�       �                    �?�S����?             3@�       �                    �?�����H�?             2@�       �       	          `ff�?z�G�z�?             $@�       �                    d@�����H�?             "@������������������������       �                     @�       �                   ht@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK�KK��ha�Bp       �t@     �x@     0r@     �b@     �p@     @V@     �A@      >@      1@              2@      >@      *@      &@      �?      $@      �?                      $@      (@      �?      (@                      �?      @      3@      �?      1@              1@      �?              @       @       @               @       @               @       @             �l@     �M@      S@      @     @R@      @      "@      @      "@      �?      @      �?              �?      @              @                       @      P@              @      @              @      @              c@      J@      2@     �@@       @      <@       @      3@              &@       @       @       @                       @              "@      0@      @      "@      @      @              @      @      @       @      @              �?       @      �?                       @              @      @             �`@      3@      3@      $@      @              *@      $@              @      *@      @      *@      �?       @      �?              �?       @              &@                      @      ]@      "@     �[@      @      [@      @     �Y@      �?      S@              ;@      �?      :@              �?      �?              �?      �?              @       @      @       @      @                       @      �?              @      @      @                      @      @      @      @               @      @       @                      @      ;@      O@      :@      D@       @     �@@       @      2@      @              @      2@              0@      @       @               @      @                      .@      2@      @      *@      �?      @      �?      �?      �?              �?      �?              @              "@              @      @      @              �?      @      �?                      @      �?      6@              4@      �?       @      �?                       @      F@      o@      9@     �l@      8@     �b@      @     @R@       @              @     @R@             �P@      @      @      @      @              @      @                      @      3@     �R@      @              ,@     �R@       @      @       @      �?              �?       @                       @      (@      R@      (@     �E@      "@      0@      @      *@      @      *@       @               @      *@               @       @      &@       @      @      �?              �?      @              �?      �?       @      �?                       @               @      �?              @      @      @                      @      @      ;@      �?      9@              3@      �?      @      �?                      @       @       @       @                       @              =@      �?      T@              R@      �?       @      �?                       @      3@      4@      ,@      @       @       @       @                       @      (@       @       @              @       @               @      @              @      0@       @              @      0@       @      0@       @       @      �?       @              @      �?       @               @      �?              �?                       @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJQY%hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK߅�h��B�0         x                    �?�Z���?�           ��@       1                    �?~�Q7:�?           �z@               	          ����?�Q����?c             d@       	       
             �?\�����?A            �[@                          �c@`���i��?             F@������������������������       �                     B@              	             �?      �?              @������������������������       �                     @������������������������       �                     �?
                          @E@�GN�z�?(            �P@                          �_@z�G�z�?             $@                          `[@�q�q�?             @������������������������       �                     �?                           �J@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           @D@      �?              L@������������������������       �                      @                           �?h�WH��?             K@                           �?�θ�?             *@������������������������       �                     @                          �q@և���X�?             @                            I@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                          �c@������?            �D@������������������������       �                     ?@                          �i@z�G�z�?             $@������������������������       �                      @������������������������       �                      @!       0       	          ����?�:pΈ��?"             I@"       -       	          ����?z�G�z�?            �A@#       $                   ``@     ��?             @@������������������������       �        
             .@%       &                    a@�t����?
             1@������������������������       �                     �?'       (                    `@      �?	             0@������������������������       �                     $@)       ,                    b@�q�q�?             @*       +                    �N@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @.       /                   �R@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@2       9                    �?X�@��l�?�            �p@3       4                   �Q@���N8�?6             U@������������������������       �                      @5       6                   `c@��Y��]�?4            �T@������������������������       �        /             S@7       8                   Pg@�q�q�?             @������������������������       �                      @������������������������       �                     @:       ]                    @L@      �?z             g@;       T       	          033�?8�Z$���?X            @`@<       Q                    @�D�d@6�?Q            �]@=       H       
             �?��ϭ�*�?N             ]@>       ?                    �?      �?             0@������������������������       �                     @@       G                   �b@�q�q�?	             (@A       B       
             �?      �?              @������������������������       �                      @C       F       	             �?�q�q�?             @D       E                   �_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @I       J                    @G@p���?B             Y@������������������������       �        !             J@K       P                   �f@ �q�q�?!             H@L       O                   @[@`Ql�R�?             �G@M       N                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �F@������������������������       �                     �?R       S                    �H@�q�q�?             @������������������������       �                      @������������������������       �                     �?U       X       	             @���!pc�?             &@V       W                    �?      �?             @������������������������       �                      @������������������������       �                      @Y       Z       	             
@؇���X�?             @������������������������       �                     @[       \                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?^       o       	          `ff�?|��?���?"             K@_       f                   �b@4�B��?            �B@`       a                    �L@d}h���?             <@������������������������       �                     @b       c                    @�8��8��?             8@������������������������       �                     4@d       e                    �?      �?             @������������������������       �                      @������������������������       �                      @g       n       	          pff�?�q�q�?             "@h       i                   �d@և���X�?             @������������������������       �                     @j       m       
             �?      �?             @k       l                   p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @p       u       	          `ff@@�0�!��?             1@q       t                    �?@4և���?             ,@r       s                    �L@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @v       w       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?y       �                    [@$��n�?�             s@z                          `n@���Q��?
             .@{       ~                   �`@�	j*D�?             *@|       }                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    �?D����?�            0r@�       �                    �?�q�����?             I@�       �                    �J@�q�q�?             B@�       �                   �a@j���� �?             1@�       �       	             �?�θ�?             *@�       �       	             �?r�q��?             (@������������������������       �                     @�       �                     I@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �O@�d�����?             3@�       �                   �`@�8��8��?	             (@�       �       	          ����?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   `f@և���X�?             @������������������������       �                     @������������������������       �                     @�       �       
             �?d}h���?             ,@�       �       	             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                    �?Ԙ-w���?�             n@�       �                   �d@<2r�Y�?�             h@�       �                   �l@�e�N�c�?�            �g@�       �       
             �?�]��?F            �Y@�       �                   �h@�x�E~�?<            @V@������������������������       �        (            �M@�       �                    �?��S�ۿ?             >@�       �       
             �?���}<S�?             7@������������������������       �                     @�       �                   p`@�KM�]�?             3@�       �                    �K@r�q��?             (@������������������������       �                     "@�       �                   pj@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �_@؇���X�?
             ,@������������������������       �                     @�       �                   p`@����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?�Ra����?;             V@������������������������       �                     3@�       �                    �R@�~t��?-            @Q@�       �       	          ����?�G�V�e�?,             Q@�       �                   Hq@ҳ�wY;�?             1@�       �                   �]@�q�q�?             "@������������������������       �                     @�       �                   0p@      �?             @�       �                   �`@      �?             @�       �                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    �?�IєX�?!            �I@�       �       	          033@�8��8��?             B@�       �                    @M@ 7���B�?             ;@������������������������       �                     6@�       �       	          `ff�?z�G�z�?             @������������������������       �                     @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          `ff
@�<ݚ�?             "@�       �                   �_@���Q��?             @�       �                   �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        	             .@������������������������       �                     �?�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �b@�q�q��?              H@�       �                   �e@���H��?             E@�       �                   �s@��(\���?             D@�       �                    �?�7��?            �C@�       �       
             �?�8��8��?             8@������������������������       �                     6@������������������������       �                      @������������������������       �        	             .@������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�        u@     �x@     Pq@     �b@     �M@     @Y@      J@      M@      �?     �E@              B@      �?      @              @      �?             �I@      .@       @       @       @      @      �?              �?      @      �?                      @              @     �H@      @               @     �H@      @      $@      @      @              @      @      @      �?              �?      @                       @     �C@       @      ?@               @       @               @       @              @     �E@      @      <@      @      ;@              .@      @      (@      �?              @      (@              $@      @       @      �?       @               @      �?              @               @      �?              �?       @                      .@     @k@      I@      T@      @               @      T@       @      S@              @       @               @      @             @a@      G@     �[@      4@     �Z@      (@     �Z@      $@       @       @      @              @       @      @      @       @               @      @      �?      @              @      �?              �?                      @     �X@       @      J@              G@       @      G@      �?      �?      �?      �?                      �?     �F@                      �?      �?       @               @      �?              @       @       @       @               @       @              �?      @              @      �?      �?      �?                      �?      <@      :@      9@      (@      6@      @              @      6@       @      4@               @       @               @       @              @      @      @      @              @      @      �?       @      �?       @                      �?      �?                       @      @      ,@      �?      *@      �?      @      �?                      @               @       @      �?       @                      �?     �N@     �n@      "@      @      "@      @      �?      @      �?                      @       @                       @      J@     �m@      :@      8@      .@      5@      $@      @      $@      @      $@       @      @              @       @               @      @                      �?              @      @      ,@      �?      &@      �?      @      �?                      @               @      @      @              @      @              &@      @      �?      @              @      �?              $@              :@     �j@      .@     @f@      ,@      f@      @     �X@       @     �U@             �M@       @      <@       @      5@              @       @      1@       @      $@              "@       @      �?       @                      �?              @              @       @      (@              @       @      @       @                      @      $@     �S@              3@      $@     �M@      "@     �M@      @      &@      @      @      @              @      @      �?      @      �?      �?      �?                      �?               @       @                       @      @      H@      @     �@@      �?      :@              6@      �?      @              @      �?      �?              �?      �?               @      @       @      @       @       @       @                       @              �?              @              .@      �?              �?      �?      �?                      �?      &@     �B@      @     �B@      @     �B@       @     �B@       @      6@              6@       @                      .@      �?               @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��fbhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK˅�h��Bh,         p                    �?�#i����?�           ��@       7       
             �?D�X%��?           �x@       0       	          pff�?h?\P��?�            �q@       +                   �a@D��2(�?r             f@                          `_@�U�����?S            ``@                           @Q@�����?)            �O@                           �?P���Q�?(             N@������������������������       �                     A@	                           �?ȵHPS!�?             :@
                          �[@�S����?             3@              	             �?      �?              @������������������������       �                     @                          @n@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     &@������������������������       �                     @������������������������       �                     @                          �k@������?*             Q@                          `f@�KM�]�?             C@                           �?���7�?             6@              
             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     *@                            L@     ��?             0@������������������������       �                     *@������������������������       �                     @       "       	             �?���Q��?             >@       !                    �?ףp=
�?             $@                            �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @#       (                    �?R���Q�?             4@$       %                   �b@�IєX�?             1@������������������������       �        
             ,@&       '                    �N@�q�q�?             @������������������������       �                      @������������������������       �                     �?)       *                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?,       /                    �H@����?�?            �F@-       .                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     C@1       6       
             �?@��!�Q�?J            @Z@2       5                     K@XB���?             =@3       4       	          033@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ;@������������������������       �        8             S@8       [       	          ����?f=UBS�?G            @]@9       X                    �?��Sݭg�?.            �S@:       ;                   �d@��X���?(            @Q@������������������������       �                      @<       =                    �?��f/w�?$            �N@������������������������       �                     *@>       K                    �L@r�qG�?             H@?       F                    �?6YE�t�?            �@@@       A                   �_@      �?              @������������������������       �                      @B       C                   0j@�q�q�?             @������������������������       �                      @D       E                    p@      �?             @������������������������       �                      @������������������������       �                      @G       H                   �b@`2U0*��?             9@������������������������       �                     5@I       J                   po@      �?             @������������������������       �                     �?������������������������       �                     @L       Q                    �?��S���?	             .@M       P                   �q@z�G�z�?             @N       O                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @R       W                    �?���Q��?             $@S       V       	          ����?�q�q�?             "@T       U                   P`@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?Y       Z                   ``@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @\       a                    �?�θ�?            �C@]       ^                    �?      �?             @������������������������       �                      @_       `                   `[@      �?              @������������������������       �                     �?������������������������       �                     �?b       i                   �`@b�h�d.�?            �A@c       d                    �?���7�?             6@������������������������       �                     $@e       h                    �?�8��8��?             (@f       g                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@j       k                    �?�n_Y�K�?
             *@������������������������       �                     @l       m                    @M@�����H�?             "@������������������������       �                     @n       o                     N@�q�q�?             @������������������������       �                     �?������������������������       �                      @q       �                    �K@,Tg�x0�?�             u@r       �       
             �?T�6|���?             j@s       x                   �Q@~h����?"             L@t       w                    �?      �?              @u       v                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @y       z                    �?�q�q�?             H@������������������������       �                     *@{       |       
             �?և���X�?            �A@������������������������       �                     @}       �                    d@     ��?             @@~       �                   0a@����X�?             5@       �                    �E@��
ц��?             *@�       �                    @C@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       	          ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?"pc�
�?             &@�       �                    @ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     �?�       �                    I@pe�D�ϣ?]             c@�       �                   �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @n@�P[1N�?[            �b@������������������������       �        7            �U@�       �                    �G@0�z��?�?$             O@�       �                   0c@XB���?             =@�       �                   �\@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@������������������������       �                    �@@�       �                   �`@     ^�?Q             `@�       �       	          pff�?�q�q�?"            �I@�       �                   @b@l��[B��?             =@�       �                   @V@��Q��?             4@�       �       
             �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?؇���X�?             ,@�       �                   @[@�q�q�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?�����H�?             "@�       �                    @r�q��?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?��2(&�?             6@�       �                   `]@և���X�?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        	             .@�       �       	          ��� @���!pc�?/            @S@�       �                   �o@r�q��?'            �P@�       �                   �a@���N8�?             E@�       �                    �?�r����?
             .@������������������������       �                     �?�       �                    �?@4և���?	             ,@�       �                   �`@ףp=
�?             $@�       �       
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     ;@�       �                   @q@      �?             8@������������������������       �                     @�       �                   �q@r�q��?             2@������������������������       �                     @�       �                    �?�θ�?             *@������������������������       �                     $@������������������������       �                     @�       �                    �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       `u@     �x@     �V@     0s@      8@     p@      7@      c@      6@     @[@      @     �L@      @     �L@              A@      @      7@      @      0@      @      @              @      @       @      @                       @              &@              @      @              0@      J@      @      A@      �?      5@      �?       @      �?                       @              *@      @      *@              *@      @              (@      2@      "@      �?      �?      �?      �?                      �?       @              @      1@      �?      0@              ,@      �?       @               @      �?               @      �?       @                      �?      �?      F@      �?      @      �?                      @              C@      �?      Z@      �?      <@      �?      �?      �?                      �?              ;@              S@     �P@      I@      M@      4@      L@      *@       @              H@      *@      *@             �A@      *@      <@      @      @      @       @               @      @               @       @       @       @                       @      8@      �?      5@              @      �?              �?      @              @       @      �?      @      �?      �?      �?                      �?              @      @      @      @      @       @      @       @                      @      @                      �?       @      @              @       @              "@      >@      @      �?       @              �?      �?              �?      �?              @      =@      �?      5@              $@      �?      &@      �?      �?      �?                      �?              $@      @       @      @              �?       @              @      �?       @      �?                       @     `o@     @U@     @f@      >@      =@      ;@      �?      @      �?      �?              �?      �?                      @      <@      4@      *@              .@      4@              @      .@      1@      @      .@      @      @      @      �?              �?      @              �?      @              @      �?                       @      "@       @      "@      �?      "@                      �?              �?     �b@      @      �?       @      �?                       @     �b@      �?     �U@             �N@      �?      <@      �?      @      �?              �?      @              6@             �@@             @R@     �K@      1@      A@      ,@      .@      *@      @      �?      @              @      �?              (@       @      @       @      �?       @      �?                       @      @               @              �?       @      �?      @              @      �?      �?              �?      �?                      @      @      3@      @      @      @      �?              �?      @                      @              .@      L@      5@     �K@      &@      D@       @      *@       @              �?      *@      �?      "@      �?      @      �?              �?      @              @              @              ;@              .@      "@              @      .@      @      @              $@      @      $@                      @      �?      $@              $@      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ$�phG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��BX)         t       
             �?"��G,�?�           ��@       !                    �?�*�@P��?            {@                           �?�G��l��?*            �O@                           �?���|���?            �@@       
                    b@����X�?
             ,@       	                     M@և���X�?             @                          `@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          �X@�KM�]�?             3@������������������������       �                     �?                          �`@�X�<ݺ?             2@                          `X@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@                           �?���Q��?             >@                          pl@$��m��?             :@              	          ����?      �?              @������������������������       �                     @������������������������       �                     @              	             �?�<ݚ�?             2@                          `^@      �?	             0@������������������������       �                     @                           �?$�q-�?             *@������������������������       �                     �?������������������������       �                     (@������������������������       �                      @                           �a@      �?             @������������������������       �                     �?������������������������       �                     @"       3                   �g@\�?A�?�            0w@#       $                    �?���f�?L             `@������������������������       �        4            @U@%       0                   �c@�Ra����?             F@&       +                    �?��p\�?            �D@'       (                   �c@�g�y��?             ?@������������������������       �                     :@)       *                    �P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?,       /                    �?z�G�z�?             $@-       .       	          ����?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @1       2                    @H@�q�q�?             @������������������������       �                     �?������������������������       �                      @4       i                   �a@d�.����?�            @n@5       D                    @K@ӏ�[��?[            @c@6       9                   @j@�?�P�a�?#             N@7       8                    �F@      �?              @������������������������       �                     @������������������������       �                     @:       A       	          033@0G���ջ?             J@;       <                    �?`���i��?             F@������������������������       �                    �B@=       @                   �]@؇���X�?             @>       ?                   @e@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @B       C                   �\@      �?              @������������������������       �                      @������������������������       �                     @E       N                   �[@�*/�8V�?8            �W@F       M       	          `ff�?��S���?             .@G       H                   �h@���|���?             &@������������������������       �                      @I       J                    l@�<ݚ�?             "@������������������������       �                     @K       L                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @O       V       	          ����?l������?0            �S@P       U                    �?�n_Y�K�?             *@Q       R       	          ����?���!pc�?             &@������������������������       �                      @S       T                   �b@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @W       h                    �?��2(&�?(            �P@X       c                   �`@�3Ea�$�?             G@Y       Z                   �h@r֛w���?             ?@������������������������       �                      @[       ^                    b@V�a�� �?             =@\       ]                   Xy@���}<S�?             7@������������������������       �                     5@������������������������       �                      @_       `                   Pb@�q�q�?             @������������������������       �                     @a       b                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?d       e                   �b@��S�ۿ?	             .@������������������������       �                     *@f       g                   `q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@j       s       	          ����?�zvܰ?1             V@k       l                    `@��2(&�?             6@������������������������       �        	             .@m       r                   @q@և���X�?             @n       o                   p`@      �?             @������������������������       �                      @p       q                     P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        $            �P@u       �                    I@DE��2{�?�            �r@v       {                    �N@؇���X�?            �A@w       x                    �M@��S�ۿ?             >@������������������������       �                     4@y       z                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @|       }                   �`@���Q��?             @������������������������       �                      @~              	          ����?�q�q�?             @������������������������       �                     �?�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��%p���?�            �p@�       �                    �?@�z�G�?4             T@�       �                   �b@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?������������������������       �        ,            �P@�       �                    �?��wv��?q             g@�       �                    �?��q縬�?b            �c@�       �                   �j@��V#�?            �E@�       �                   pc@�n_Y�K�?             *@������������������������       �                     @������������������������       �                      @�       �                   �b@z�G�z�?             >@�       �       	          ����?PN��T'�?             ;@�       �                   �q@ףp=
�?             4@������������������������       �        	             .@�       �                   �_@���Q��?             @������������������������       �                      @������������������������       �                     @�       �       	          ����?����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �E@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @[@,Z0R�?H             ]@�       �                    �G@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �g@@-�_ .�?F            �[@�       �                   �c@���7�?E            �[@�       �                    @L@Pa�	�??            �X@������������������������       �        2            @S@�       �                   �a@��2(&�?             6@������������������������       �                     (@�       �                   �a@�z�G��?             $@������������������������       �                      @�       �                    b@      �?              @�       �       	             �?�q�q�?             @�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �p@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @������������������������       �                     �?�       �                   @`@�n_Y�K�?             :@������������������������       �                     @�       �                    �?      �?             4@�       �                    �?r�q��?             (@�       �       	             �?�<ݚ�?             "@�       �                   `k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       @s@     �z@      R@     �v@     �@@      >@      5@      (@      @      $@      @      @      �?      @              @      �?              @                      @      1@       @              �?      1@      �?      @      �?              �?      @              $@              (@      2@      "@      1@      @      @      @                      @      @      ,@      @      (@      @              �?      (@      �?                      (@               @      @      �?              �?      @             �C@     �t@      @      _@             @U@      @     �C@      @      C@      �?      >@              :@      �?      @              @      �?               @       @       @       @       @                       @              @       @      �?              �?       @              A@      j@      ?@     �^@      @     �J@      @      @      @                      @      @     �H@      �?     �E@             �B@      �?      @      �?       @      �?                       @              @       @      @       @                      @      8@     �Q@      @       @      @      @               @      @       @      @              �?       @               @      �?                      @      1@      O@       @      @       @      @               @       @      �?       @                      �?               @      "@     �L@      "@     �B@       @      7@       @              @      7@       @      5@              5@       @              @       @      @              �?       @               @      �?              �?      ,@              *@      �?      �?      �?                      �?              4@      @     @U@      @      3@              .@      @      @      @      �?       @              �?      �?      �?                      �?              @             �P@     �m@      P@      @      >@       @      <@              4@       @       @       @                       @      @       @       @              �?       @              �?      �?      �?      �?                      �?     �l@      A@     �S@      �?      (@      �?      (@                      �?     �P@              c@     �@@      a@      7@      =@      ,@      @       @      @                       @      8@      @      7@      @      2@       @      .@              @       @               @      @              @       @               @      @              �?       @               @      �?             �Z@      "@       @      @              @       @             @Z@      @     @Z@      @      X@      @     @S@              3@      @      (@              @      @               @      @      �?       @      �?      �?      �?      �?                      �?      �?              @              "@       @      "@                       @              �?      0@      $@      @              $@      $@       @      $@       @      @       @      �?              �?       @                      @              @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJW:+LhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKǅ�h��B�+         J                   �`@�#i����?�           ��@       5                    �?p�L���?�            `s@       &       
             �?H0sE�d�?�             l@                          �`@�0p<���?             h@                          �Q@�*/�8V�?A            �W@������������������������       �                     �?              	          033@��a�n`�?@            @W@       	                   �h@���}<S�??             W@������������������������       �                     C@
              	          ����?PN��T'�?"             K@                            L@ �o_��?             9@                          �r@�8��8��?             (@������������������������       �                     $@                          @_@      �?              @������������������������       �                     �?������������������������       �                     �?                            P@��
ц��?             *@                          �\@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          `_@XB���?             =@������������������������       �                     4@                           �?�����H�?             "@                          j@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?       %       	          ����?`�LVXz�?>            �X@                            �?@4և���?
             ,@������������������������       �                     @!       $                    �L@�����H�?             "@"       #                    Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        4            @U@'       ,                   �]@     ��?             @@(       +                   Pg@�q�q�?             (@)       *       	          ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @-       .                   �_@      �?             4@������������������������       �                     &@/       4                    �?X�<ݚ�?             "@0       3       	          @33�?r�q��?             @1       2                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @6       A       
             �?k�q��?7            @U@7       <                    �?D>�Q�?"             J@8       ;                     P@      �?             (@9       :                    @�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @=       >                     Q@��(\���?             D@������������������������       �                     ?@?       @                   `_@�q�q�?             "@������������������������       �                     @������������������������       �                     @B       G                    �?�C��2(�?            �@@C       D                    @XB���?             =@������������������������       �                     ;@E       F                    @N@      �?              @������������������������       �                     �?������������������������       �                     �?H       I                    �?      �?             @������������������������       �                      @������������������������       �                      @K       V                   @E@������?
           �z@L       M                    �?z�G�z�?             >@������������������������       �                     0@N       U                   �d@և���X�?
             ,@O       T                    @      �?             (@P       S                   �^@�q�q�?             "@Q       R                   �a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @W       �                    �?�O&��<�?�            �x@X       y                    �?����p�?V             a@Y       x       	          `ff@؀�:M�?/            �R@Z       m                   `@�q�q�?,            @Q@[       h                   �^@l��[B��?             =@\       e                   �c@�ՙ/�?             5@]       `                   @l@��
ц��?	             *@^       _                     K@r�q��?             @������������������������       �                     @������������������������       �                     �?a       d                   0q@����X�?             @b       c       	          ����?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?f       g                     E@      �?              @������������������������       �                     �?������������������������       �                     @i       l                   �d@      �?              @j       k                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @n       u       
             �?z�G�z�?             D@o       p       	          ����?      �?             (@������������������������       �                     @q       r       	          @33�?�q�q�?             "@������������������������       �                     @s       t                    �?      �?             @������������������������       �                     �?������������������������       �                     @v       w                    �M@@4և���?             <@������������������������       �                     :@������������������������       �                      @������������������������       �                     @z       �                   `\@�z�6�?'             O@{       |                     E@���Q��?             $@������������������������       �                     @}       �                   �a@և���X�?             @~              	             �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                   �s@D>�Q�?"             J@�       �                   �d@�����H�?            �F@�       �                   �b@�C��2(�?             F@�       �                    �?�X�<ݺ?             B@�       �                   8p@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     <@�       �                    @I@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    c@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �`@�1iJ�?�             p@�       �                    @L@�s�c���?d            @c@�       �       
             �?�<_���?X             a@�       �                   @^@�q�q�?             >@�       �                   �a@      �?             4@������������������������       �                     @�       �                    @j���� �?             1@�       �                    @G@����X�?
             ,@�       �       	              @z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     $@�       �                    �?���1��?D            �Z@������������������������       �                    �A@�       �                    c@�k~X��?+             R@�       �                    �?��?^�k�?            �A@������������������������       �                     (@�       �                   �b@�nkK�?             7@������������������������       �        
             6@������������������������       �                     �?������������������������       �                    �B@�       �                    �?�t����?             1@�       �       	              @X�Cc�?
             ,@�       �                    �L@"pc�
�?             &@������������������������       �                     �?�       �                    �M@ףp=
�?             $@�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       
             �?R�}e�.�?:             Z@�       �                   �b@��Q��?             D@�       �                   e@П[;U��?             =@������������������������       �                     @�       �                    �?�q�����?             9@�       �                   �q@     ��?             0@������������������������       �                     *@������������������������       �                     @������������������������       �                     "@�       �                   �l@�C��2(�?             &@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   �t@      �?'             P@������������������������       �        %            �M@�       �                   �u@���Q��?             @������������������������       �                      @������������������������       �                     @�t�b�i     h�h*h-K ��h/��R�(KK�KK��ha�Bp       `u@     �x@     �O@     �n@      8@      i@      &@     �f@      $@      U@      �?              "@      U@       @      U@              C@       @      G@      @      2@      �?      &@              $@      �?      �?      �?                      �?      @      @      @      �?              �?      @                      @      �?      <@              4@      �?       @      �?      @      �?                      @              @      �?              �?     �X@      �?      *@              @      �?       @      �?       @               @      �?                      @             @U@      *@      3@       @      @      �?      @      �?                      @      @              @      .@              &@      @      @      @      �?       @      �?       @                      �?      @                      @     �C@      G@      "@     �E@      @      @      @      @              @      @              @              @     �B@              ?@      @      @              @      @              >@      @      <@      �?      ;@              �?      �?              �?      �?               @       @       @                       @     pq@      b@      @      8@              0@      @       @      @      @      @      @      �?      @      �?                      @      @                      @               @     q@     @^@     �M@     @S@      G@      <@      G@      7@      ,@      .@      *@       @      @      @      �?      @              @      �?              @       @      @      �?      @                      �?              �?      @      �?              �?      @              �?      @      �?       @      �?                       @              @      @@       @      @      @              @      @      @      @              �?      @      �?                      @      :@       @      :@                       @              @      *@     �H@      @      @              @      @      @      @       @      @                       @              �?      "@     �E@      @      D@      @      D@       @      A@       @      @       @                      @              <@       @      @       @                      @      �?              @      @              @      @             �j@      F@     @a@      0@     �_@      &@      4@      $@      $@      $@              @      $@      @      $@      @       @       @       @                       @       @       @       @                       @              @      $@             �Z@      �?     �A@             �Q@      �?      A@      �?      (@              6@      �?      6@                      �?     �B@              (@      @      "@      @      "@       @              �?      "@      �?      @      �?      @                      �?      @                      @      @              S@      <@      ,@      :@      *@      0@              @      *@      (@      *@      @      *@                      @              "@      �?      $@      �?      �?      �?                      �?              "@      O@       @     �M@              @       @               @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJF<KdhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B�'         b       
             �?�#i����?�           ��@       I                   �b@L�~m��?           �x@       (                    �?�Zl�i��?�            @t@                           b@���D�?�            �l@������������������������       �        *             O@       %                    �Q@�8��8��?p             e@       $                    �?�u�w�u�?m            `d@              	          ����?����y7�?V            @_@	                           �?�%^�?            �E@
              	          ����?�θ�?            �C@������������������������       �        	             3@                           �?�G�z��?             4@                          �`@�<ݚ�?             "@������������������������       �                     @                           �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?���|���?
             &@                          `c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?                           @K@      �?             @������������������������       �                      @              	             �?      �?             @������������������������       �                     @������������������������       �                     �?                          @^@      �?             @������������������������       �                      @������������������������       �                      @       #                   �\@����ȫ�?:            �T@       "                   �`@      �?              @        !                    �K@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        6            �R@������������������������       �                     C@&       '                   �]@���Q��?             @������������������������       �                     @������������������������       �                      @)       2                    �?��k=.��?;            �W@*       +       	             �?���Q��?
             .@������������������������       �                     @,       1                    @ףp=
�?             $@-       0       	          ����?r�q��?             @.       /                   �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @3       F                   �e@���!���?1            �S@4       5                   �]@h��@D��?.            �Q@������������������������       �                     9@6       E       	          ����?*
;&���?!             G@7       8                   �\@b�2�tk�?             2@������������������������       �                     @9       :                   �_@��S���?             .@������������������������       �                     @;       <       
             �?�q�q�?             (@������������������������       �                     �?=       >       	          ����?���!pc�?
             &@������������������������       �                     @?       @                     M@      �?             @������������������������       �                      @A       D                    �?      �?             @B       C                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     <@G       H                    �?      �?              @������������������������       �                      @������������������������       �                     @J       Q                    �?)O���?-             R@K       P                    �M@�+e�X�?             9@L       O                   �`@���Q��?	             .@M       N                   �r@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @������������������������       �                     $@R       a       	             @(���@��?            �G@S       T                    �F@���N8�?             E@������������������������       �                     &@U       V                   @J@�4�����?             ?@������������������������       �                     @W       \                    �?      �?             <@X       Y       	          033�?�}�+r��?             3@������������������������       �        	             0@Z       [                   �m@�q�q�?             @������������������������       �                      @������������������������       �                     �?]       `                    �?�q�q�?             "@^       _                   `b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @c       j                    �?4>���?�             u@d       i       	          `ff�?���N8�?6             U@e       f                   d@��Y��]�?5            �T@������������������������       �        !             H@g       h                   0d@�IєX�?             A@������������������������       �                      @������������������������       �                     @@������������������������       �                      @k       �                    �?�U���?�            �o@l       �                    �?Zz�����?5            @U@m       v                    @F@�w��#��?!             I@n       u                   �_@�q�q�?             (@o       t                   �a@z�G�z�?             $@p       q                   �\@�q�q�?             @������������������������       �                     �?r       s                   @]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @w       x                    X@�I�w�"�?             C@������������������������       �                     @y       �                    b@b�h�d.�?            �A@z       }                   �c@�r����?             >@{       |                   @E@ �q�q�?             8@������������������������       �                     �?������������������������       �                     7@~       �                   �`@      �?             @       �                     H@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �j@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �`@��R[s�?            �A@�       �                   �`@���Q��?
             .@�       �                    �?�	j*D�?	             *@�       �       	             �?և���X�?             @������������������������       �                      @�       �                    �?���Q��?             @������������������������       �                      @�       �                    S@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �k@R���Q�?
             4@�       �                   �d@�q�q�?             "@�       �                   pj@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                   �t@��C[���?c             e@�       �       	             @�5U��K�?b            �d@�       �                    @�>����?`            @d@�       �                    �?@-�_ .�?Y            �b@�       �                    �?���tcH�?K            @^@�       �                    @L@ �Jj�G�?'            �K@������������������������       �                     �G@�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     @�       �                   @[@�FVQ&�?$            �P@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        "             N@�       �                    �Q@�����H�?             ;@������������������������       �                     8@������������������������       �                     @�       �                   �b@����X�?             ,@�       �                   @`@ףp=
�?             $@�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h*h-K ��h/��R�(KK�KK��ha�BP       `u@     �x@     �Q@     `t@      @@     @r@      ,@      k@              O@      ,@     @c@      (@     �b@      (@     @\@      &@      @@      "@      >@              3@      "@      &@       @      @              @       @      �?       @                      �?      @      @      @      �?      @                      �?      @      @               @      @      �?      @                      �?       @       @               @       @              �?     @T@      �?      @      �?      @              @      �?                      @             �R@              C@       @      @              @       @              2@      S@      "@      @              @      "@      �?      @      �?       @      �?              �?       @              @              @              "@     �Q@      @      P@              9@      @     �C@      @      &@              @      @       @      @              @       @      �?              @       @              @      @      @               @      @      �?      �?      �?      �?                      �?       @                      <@       @      @       @                      @      C@      A@      @      3@      @      "@      �?      "@              "@      �?              @                      $@      @@      .@      @@      $@      &@              5@      $@              @      5@      @      2@      �?      0@               @      �?       @                      �?      @      @      @       @      @                       @              @              @      q@     �P@      T@      @      T@       @      H@              @@       @               @      @@                       @      h@      O@      E@     �E@     �@@      1@      @       @       @       @       @      �?      �?              �?      �?      �?                      �?              @       @              =@      "@              @      =@      @      :@      @      7@      �?              �?      7@              @      @      �?      @      �?                      @       @              @       @               @      @              "@      :@      @      "@      @      "@      @      @       @               @      @               @       @      �?       @                      �?              @       @              @      1@      @      @      �?      @              @      �?               @                      &@     �b@      3@     �b@      0@     �b@      (@     �a@       @      ]@      @      K@      �?     �G@              @      �?              �?      @              O@      @       @      @              @       @              N@              8@      @      8@                      @      $@      @      "@      �?      �?      �?      �?                      �?       @              �?      @              @      �?                      @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJؽ�hG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B�)         h                    �?�/�$�y�?�           ��@       9       
             �?@�0�!��?�            px@       6                    �R@P�#L5ھ?�            pr@                           �?P����?�            @r@                          �`@"pc�
�?             F@                           �?8����?             7@������������������������       �                     @                           �?z�G�z�?             4@	                          a@�q�q�?             (@
                           @H@�q�q�?             @������������������������       �                     �?              	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                          `c@���N8�?             5@                           �I@$�q-�?             *@                            F@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                          �h@��d�?�             o@������������������������       �        @            @Y@                          @Z@��<D�m�?]            `b@������������������������       �                     �?                          0i@F��}��?\            @b@������������������������       �                     �?       1       	          033@�2c�$��?[             b@       &                    ]@`J����?N            �^@        %                   �e@؇���X�?             ,@!       "                   �`@$�q-�?             *@������������������������       �                     "@#       $       	             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?'       *       
             �?����q�?F            @[@(       )                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @+       ,                   @c@�K}��?@            �Y@������������������������       �        <             X@-       .       	             �?r�q��?             @������������������������       �                      @/       0                   �o@      �?             @������������������������       �                     �?������������������������       �                     @2       5       	          ���@��2(&�?             6@3       4                    �J@      �?             (@������������������������       �                     @������������������������       �                     "@������������������������       �                     $@7       8       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?:       G                   �]@�q���?C             X@;       F       	          833�?�q�q�?             8@<       A                   g@��
ц��?
             *@=       >                    @D@z�G�z�?             @������������������������       �                      @?       @                   �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @B       C                   �[@      �?              @������������������������       �                     @D       E                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@H       [       	          ����?P��E��?3             R@I       J                   `c@:�&���?            �C@������������������������       �                     0@K       Z                   �b@8����?             7@L       M                    �?z�G�z�?             4@������������������������       �                      @N       U                    �?�q�q�?	             (@O       P                   Pe@�<ݚ�?             "@������������������������       �                     @Q       T                    �?      �?             @R       S                    �J@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?V       W                    �E@�q�q�?             @������������������������       �                     �?X       Y                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @\       ]                    `@�q�q�?            �@@������������������������       �                     &@^       c                    �?      �?             6@_       `                   �d@      �?              @������������������������       �                     @a       b                    �G@      �?              @������������������������       �                     �?������������������������       �                     �?d       e                     L@����X�?	             ,@������������������������       �                     @f       g                    @N@և���X�?             @������������������������       �                     @������������������������       �                     @i       �       
             �?0�����?�            pu@j       �                    �?�*;L�?N             ^@k       �                   0r@rr�J��?0            �R@l       u       	          ����?.Lj���?,             Q@m       p                    �?�t����?	             1@n       o                     H@�q�q�?             @������������������������       �                      @������������������������       �                     �?q       r                   �m@@4և���?             ,@������������������������       �                     &@s       t                   �\@�q�q�?             @������������������������       �                      @������������������������       �                     �?v       �                   �o@j���� �?#            �I@w       �       	          ��� @�\��N��?             C@x                           `@ �o_��?             9@y       z                    �K@�eP*L��?             &@������������������������       �                     @{       ~                    �?      �?              @|       }                   �_@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                   0a@؇���X�?             ,@������������������������       �                     "@�       �                   pc@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   @n@8�Z$���?             *@�       �       
             �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?�       �                    �K@$�q-�?	             *@�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     @�       �                   �`@�㙢�c�?             G@�       �       
             �?      �?             @@������������������������       �                     @�       �                   P`@XB���?             =@�       �       	             �?�����H�?             "@������������������������       �                     @�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@�       �                    \@      �?
             ,@������������������������       �                     �?�       �                    �I@��
ц��?	             *@�       �                    �D@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     @������������������������       �                     @�       �                    @h�qVhԳ?�            �k@�       �       	          ���@��.N"Ҭ?|            �i@�       �                   @g@ R�,3��?z            �i@�       �       	            �? ��ʻ��?y            �i@�       �                   �c@���ib#�?f            �e@�       �                   �t@@�K�҈?_            �d@������������������������       �        ]             d@�       �                   y@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   `_@�C��2(�?             &@�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   �a@XB���?             =@�       �                   @a@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     1@������������������������       �                     �?������������������������       �                      @�       �                   Pp@     ��?	             0@�       �                   0i@@4և���?             ,@������������������������       �                     "@�       �                   �j@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�        t@     �y@     @Q@      t@      3@     @q@      1@     0q@       @      B@      @      0@      @              @      0@      @       @      @       @              �?      @      �?      @                      �?              @               @      �?      4@      �?      (@      �?      @              @      �?                       @               @      "@     �m@             @Y@      "@     @a@      �?               @     @a@      �?              @     @a@      @     �]@       @      (@      �?      (@              "@      �?      @              @      �?              �?               @     �Z@      �?      @      �?                      @      �?     @Y@              X@      �?      @               @      �?      @      �?                      @      @      3@      @      "@      @                      "@              $@       @      �?       @                      �?      I@      G@      @      1@      @      @      �?      @               @      �?       @      �?                       @      @       @      @              �?       @               @      �?                      &@     �E@      =@      @@      @      0@              0@      @      0@      @       @               @      @      @       @      @               @       @      �?       @      �?                       @      �?              �?       @              �?      �?      �?              �?      �?                      @      &@      6@              &@      &@      &@      @      �?      @              �?      �?      �?                      �?      @      $@              @      @      @      @                      @     `o@      W@     �B@     �T@      =@     �F@      7@     �F@       @      .@      �?       @               @      �?              �?      *@              &@      �?       @               @      �?              5@      >@      4@      2@      2@      @      @      @              @      @       @      @       @      @                       @       @              (@       @      "@              @       @      @                       @       @      &@      �?      &@      �?                      &@      �?              �?      (@      �?       @      �?                       @              $@      @               @      C@      �?      ?@              @      �?      <@      �?       @              @      �?      �?              �?      �?                      4@      @      @      �?              @      @      �?      @      �?                      @      @      @      @                      @     �j@      "@      i@      @      i@      @      i@      @     �e@       @     `d@      �?      d@               @      �?              �?       @              $@      �?      �?      �?              �?      �?              "@              <@      �?      &@      �?      &@                      �?      1@                      �?               @      *@      @      *@      �?      "@              @      �?              �?      @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJX��vhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B�$         X       
             �?���
%�?�           ��@       3                    �? ��7E��?           �z@              	          ����?�Kǔ�{�?f            `d@                           @E@ pƵHP�?              J@                          pe@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     F@	       &                   �`@��_����?F            �[@
                           \@     8�?'             P@                           �M@����X�?             @������������������������       �                      @������������������������       �                     @                          �Z@�^���U�?"            �L@������������������������       �                     "@                          k@r�qG�?             H@              	          `ff@�����?             5@                          �^@�X�<ݺ?             2@              
             �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@                          �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?�5��?             ;@              	          ����?؇���X�?             @������������������������       �                     �?������������������������       �                     @       !                    m@      �?
             4@                            �?և���X�?             @������������������������       �                     @������������������������       �                     @"       #                    �?$�q-�?             *@������������������������       �                     $@$       %                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @'       2                    �R@dP-���?            �G@(       +                    a@���.�6�?             G@)       *                    �?      �?              @������������������������       �                      @������������������������       �                     @,       1       
             �?P�Lt�<�?             C@-       0                    ]@�����H�?             "@.       /                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     =@������������������������       �                     �?4       =                    �?�iyw	
�?�            �p@5       <                    �J@��a�n`�?             ?@6       7                   h@���|���?             &@������������������������       �                     @8       9       	          ����?      �?              @������������������������       �                     @:       ;                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             4@>       O       	          ����?8�M'��?�            �m@?       @                   `h@�C��2(�?3            @S@������������������������       �                    �C@A       B       	          ����?>A�F<�?             C@������������������������       �                     .@C       D                    �?8����?             7@������������������������       �                      @E       F       	             �?�q�q�?             5@������������������������       �                      @G       H                   �[@�d�����?             3@������������������������       �                     �?I       J                    �?�<ݚ�?             2@������������������������       �        	             *@K       N                     M@z�G�z�?             @L       M                   m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @P       U                   Ps@�(\����?c             d@Q       T                   0c@PL��V�?\            �b@R       S                   �Z@�-�|�?[            `b@������������������������       �                      @������������������������       �        Y             b@������������������������       �                     �?V       W       
             �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@Y       �                    �?�˱��H�?�            �r@Z       k                    �?fK!���?6            �V@[       `                   @\@����"�?             =@\       _       	          ����?�����H�?             "@]       ^                   �_@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @a       h       	          033�?      �?             4@b       e                    �L@     ��?
             0@c       d                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @f       g                   f@r�q��?             @������������������������       �                     @������������������������       �                     �?i       j                   �b@      �?             @������������������������       �                     @������������������������       �                     �?l              	             �?�P�*�?%             O@m       x                    �?�GN�z�?             F@n       s                    �?<���D�?            �@@o       p                   �e@XB���?             =@������������������������       �                     ;@q       r                    @C@      �?              @������������������������       �                     �?������������������������       �                     �?t       w                    �?      �?             @u       v                    ]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @y       z                    �?�eP*L��?             &@������������������������       �                     @{       |                    �M@      �?              @������������������������       �                     @}       ~                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          `ff�?�����H�?             2@������������������������       �        	             0@������������������������       �                      @�       �                   �g@ �h�7W�?�            �j@�       �                   p`@P�S�L�?�            `j@�       �                    @G@������?X             b@������������������������       �        (            �P@�       �       	             @�7��?0            �S@�       �                    �G@`<)�+�?/            @S@������������������������       �                      @�       �                    �?�}��L�?.            �R@������������������������       �                     >@�       �                   (p@����?�?            �F@������������������������       �                     A@�       �                    @L@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     �?�       �       	          ����?pH����?4            �P@�       �                    @ ��WV�?)             J@�       �                    �?@��8��?%             H@������������������������       �        
             *@�       �                    �?��?^�k�?            �A@�       �                   �a@h�����?             <@�       �                   xt@      �?             0@������������������������       �                     .@������������������������       �                     �?������������������������       �        	             (@������������������������       �                     @�       �                    @N@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �l@�q�q�?             .@�       �                   pb@X�<ݚ�?             "@�       �                    d@����X�?             @�       �                    �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�
       0s@     �z@      N@     0w@      E@     @^@      �?     �I@      �?      @              @      �?                      F@     �D@     �Q@     �B@      ;@       @      @       @                      @     �A@      6@              "@     �A@      *@      3@       @      1@      �?      @      �?              �?      @              $@               @      �?       @                      �?      0@      &@      �?      @      �?                      @      .@      @      @      @              @      @              (@      �?      $@               @      �?              �?       @              @     �E@      @     �E@       @      @       @                      @      �?     �B@      �?       @      �?      �?      �?                      �?              @              =@      �?              2@     @o@      @      8@      @      @      @              @      @      @              �?      @              @      �?                      4@      &@     @l@      @     �Q@             �C@      @      ?@              .@      @      0@               @      @      ,@       @              @      ,@      �?              @      ,@              *@      @      �?      �?      �?      �?                      �?      @              @     �c@      @      b@       @      b@       @                      b@      �?              �?      &@      �?                      &@     �n@      L@     �G@      F@      &@      2@      �?       @      �?      @      �?                      @              @      $@      $@      "@      @       @       @       @                       @      �?      @              @      �?              �?      @              @      �?              B@      :@      A@      $@      =@      @      <@      �?      ;@              �?      �?      �?                      �?      �?      @      �?      �?      �?                      �?               @      @      @      @               @      @              @       @      �?       @                      �?       @      0@              0@       @              i@      (@      i@      &@     �a@      @     �P@             �R@      @     �R@      @               @     �R@      �?      >@              F@      �?      A@              $@      �?      $@                      �?              �?      N@      @      I@       @     �G@      �?      *@              A@      �?      ;@      �?      .@      �?      .@                      �?      (@              @              @      �?              �?      @              $@      @      @      @       @      @       @      �?       @                      �?              @       @              @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���EhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKم�h��Bx/         ^       	          033�?�r,��?�           ��@       +       
             �?H;N	�	�?�             x@       
                   �g@�&�5y�?J             _@                           �?`���i��?             F@������������������������       �                    �A@                          `]@�����H�?             "@������������������������       �                     @       	                     @�q�q�?             @������������������������       �                     �?������������������������       �                      @       $                    �?��Q��?.             T@                           @D@~h����?              L@������������������������       �                     "@              	          ����?֭��F?�?            �G@              
             �?���N8�?             5@������������������������       �                      @                           @E@�S����?             3@������������������������       �                     �?                           @P@�����H�?             2@                           �H@�IєX�?             1@                            H@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?                          �b@$�q-�?             :@������������������������       �                     $@              	          833�?      �?             0@������������������������       �                     @              	          ����?z�G�z�?             $@������������������������       �                     �?        #                     J@�����H�?             "@!       "                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @%       (                     H@r�q��?             8@&       '                   @q@�q�q�?             @������������������������       �                      @������������������������       �                     �?)       *                   �Z@�����?             5@������������������������       �                      @������������������������       �                     3@,       ;                   @E@8Ӈ���?�            `p@-       :       	          hff�?8�A�0��?             6@.       9                    d@������?
             1@/       8                   �c@�r����?	             .@0       1                   �`@@4և���?             ,@������������������������       �                     "@2       3                    �?z�G�z�?             @������������������������       �                     �?4       5                   �]@      �?             @������������������������       �                      @6       7                   0a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @<       O                    �?��(\���?�             n@=       D                    c@r�qG�?              H@>       ?                   �j@�t����?             1@������������������������       �                     �?@       A                    q@      �?
             0@������������������������       �                     *@B       C                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?E       N                   �b@f���M�?             ?@F       M                   �_@������?             ;@G       H                    �?      �?	             ,@������������������������       �                     @I       J                   `\@�<ݚ�?             "@������������������������       �                     @K       L                   �^@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        
             *@������������������������       �                     @P       [                   �t@��8����?}             h@Q       R                   d@�~��?y            �f@������������������������       �        L             \@S       V                   Pd@����Q8�?-            �Q@T       U                   �_@      �?             @������������������������       �                     @������������������������       �                     @W       Z                    �? ����?)            @P@X       Y                    k@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        &            �N@\       ]                   u@�����H�?             "@������������������������       �                     �?������������������������       �                      @_       �                   �b@д>��C�?�            �u@`       �                   P`@܍�l�p�?�             r@a       j                    �?�P��G7�?Q            @]@b       c                   �Z@և���X�?             ,@������������������������       �                     @d       i                     K@z�G�z�?             $@e       f                    �?���Q��?             @������������������������       �                      @g       h                    @I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @k       �                    �?�	��)��?I            �Y@l       �       	          ��� @x!'ǯ�?8            �R@m       n                    V@x��}�?(            �K@������������������������       �                     �?o       |                    @L@�<ݚ�?'             K@p       y                    �?ܷ��?��?             =@q       r                    �?�nkK�?             7@������������������������       �                     @s       x                   �[@P���Q�?             4@t       w                    b@r�q��?             @u       v                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@z       {                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @}       �                   �^@��H�}�?             9@~       �                    @z�G�z�?             .@       �                    �L@؇���X�?
             ,@������������������������       �                     �?�       �       	             �?$�q-�?	             *@������������������������       �                     &@�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   @`@���Q��?             $@�       �                   `]@      �?              @�       �                   `Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   �Z@�KM�]�?             3@�       �                   d@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�IєX�?             1@������������������������       �                     .@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     =@�       �                    �?Pt�nٔ�?e            �e@�       �                   �s@ȵHPS!�?             :@�       �                    @HP�s��?             9@������������������������       �                     3@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �       
             �?��<�Ұ?V            `b@�       �                    �?`���i��?P            �`@�       �                    �?���1��??            �Z@�       �                    �?$�q-�?             *@������������������������       �                     @�       �                    �H@؇���X�?             @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        8            �W@�       �                   �`@HP�s��?             9@������������������������       �                     3@�       �                    �?�q�q�?             @�       �       	             @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    S@�r����?             .@�       �                    �L@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    \@      �?&             M@������������������������       �                     @�       �                    �L@�>���?#             K@�       �                    �?<ݚ)�?             B@�       �                   `c@d}h���?             <@�       �                    �?8�Z$���?             :@�       �                    �?և���X�?             @�       �                   �l@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?�}�+r��?             3@�       �       	          ���@�8��8��?	             (@������������������������       �                     "@�       �                    @B@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �       
             �?      �?              @������������������������       �                     @������������������������       �                     @�       �                    �P@�<ݚ�?             2@�       �                    �?@4և���?	             ,@�       �                    �N@؇���X�?             @������������������������       �                      @�       �       	          ����?z�G�z�?             @�       �                   ps@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�t�bh�h*h-K ��h/��R�(KK�KK��ha�B�       �t@     Py@     �p@     @]@      A@     �V@      �?     �E@             �A@      �?       @              @      �?       @      �?                       @     �@@     �G@      =@      ;@              "@      =@      2@      @      0@       @              @      0@      �?               @      0@      �?      0@      �?      @              @      �?                      (@      �?              8@       @      $@              ,@       @      @               @       @              �?       @      �?       @      �?       @                      �?      @              @      4@       @      �?       @                      �?       @      3@       @                      3@     `m@      ;@      *@      "@      *@      @      *@       @      *@      �?      "@              @      �?      �?              @      �?       @              �?      �?              �?      �?                      �?               @              @     �k@      2@     �A@      *@      .@       @              �?      .@      �?      *@               @      �?       @                      �?      4@      &@      4@      @      @      @      @               @      @              @       @      @       @                      @      *@                      @     `g@      @     `f@      @      \@             �P@      @      @      @      @                      @      P@      �?      @      �?      @                      �?     �N@               @      �?              �?       @              N@      r@      ?@     0p@      7@     �W@       @      @              @       @       @      @       @       @              �?       @      �?                       @      @              .@      V@      .@     �M@      *@      E@      �?              (@      E@      @      :@      �?      6@              @      �?      3@      �?      @      �?       @               @      �?                      @              ,@       @      @       @                      @      "@      0@      @      (@       @      (@      �?              �?      (@              &@      �?      �?      �?                      �?      �?              @      @      @       @      �?       @      �?                       @      @                       @       @      1@      �?      �?              �?      �?              �?      0@              .@      �?      �?      �?                      �?              =@       @     �d@      @      7@       @      7@              3@       @      @       @                      @      �?              @     �a@      @      `@      �?     �Z@      �?      (@              @      �?      @      �?      �?      �?                      �?              @             �W@       @      7@              3@       @      @       @      �?       @                      �?              @       @      *@       @      @              @       @                      @      =@      =@              @      =@      9@      9@      &@      6@      @      6@      @      @      @      @      �?              �?      @                       @      2@      �?      &@      �?      "@               @      �?              �?       @              @                       @      @      @      @                      @      @      ,@      �?      *@      �?      @               @      �?      @      �?      �?              �?      �?                      @              @      @      �?      @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ:9)bhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KK���h��B�(         x                    �?T8���?�           ��@       _                    �?�yZ����?           �z@       L       	          033�?���X�K�?�            �v@       )       
             �?����j��?�            �s@                          `]@�ހ��?:            �W@������������������������       �                     6@                           �?r�q��?.             R@                          �c@���}<S�?             7@	       
                   �[@z�G�z�?	             $@������������������������       �                     �?                           �?�����H�?             "@������������������������       �                     @                           c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@              	          833�?f�Sc��?            �H@              
             �?V�a�� �?             =@������������������������       �                     @                            E@ȵHPS!�?             :@                           �C@�θ�?             *@������������������������       �                     "@                          �b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@       $       	          ����?���Q��?             4@                          �_@8�Z$���?	             *@                          �^@      �?              @������������������������       �                     �?������������������������       �                     �?        !                   �c@�C��2(�?             &@������������������������       �                      @"       #                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @%       (                     F@؇���X�?             @&       '                   Pp@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @*       K                   �g@��X��?�             l@+       B                   �b@���l��?�            �k@,       -                    �?��d5z�?�            `i@������������������������       �        $             K@.       1                    X@l������?\            �b@/       0                   �[@�q�q�?             @������������������������       �                      @������������������������       �                     @2       A                    @d�;�s��?Y            �a@3       <                    _@���.�d�?X            �a@4       7                    �?�J�4�?#             I@5       6                    ]@      �?              @������������������������       �                     @������������������������       �                     @8       ;                   �a@�����?             E@9       :                   @^@�	j*D�?
             *@������������������������       �                     "@������������������������       �                     @������������������������       �                     =@=       >                    �?�����?5             W@������������������������       �        "            �L@?       @                   Pt@��?^�k�?            �A@������������������������       �                     A@������������������������       �                     �?������������������������       �                     �?C       F                    @E@���y4F�?             3@D       E                   �a@      �?             @������������������������       �                      @������������������������       �                      @G       H                    @�r����?
             .@������������������������       �                     (@I       J                    ^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @M       Z                   �d@0,Tg��?             E@N       U                     H@@�0�!��?             A@O       T                   �a@      �?              @P       Q                    �?z�G�z�?             @������������������������       �                     @R       S                   @a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @V       W                    @$�q-�?             :@������������������������       �                     6@X       Y                   �a@      �?             @������������������������       �                      @������������������������       �                      @[       \       	             @      �?              @������������������������       �                     @]       ^       
             �?���Q��?             @������������������������       �                      @������������������������       �                     @`       o       
             �?=��T�?1            �Q@a       f                    �?4?,R��?             B@b       e                   `R@ ��WV�?             :@c       d                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     8@g       l                    @O@���Q��?             $@h       i       	             �?r�q��?             @������������������������       �                     @j       k                    \@      �?              @������������������������       �                     �?������������������������       �                     �?m       n       	          ����?      �?             @������������������������       �                     �?������������������������       �                     @p       u                    �?ҳ�wY;�?             A@q       r                     G@r�q��?	             (@������������������������       �                     @s       t                    ]@����X�?             @������������������������       �                     @������������������������       �                      @v       w       	          hff @�C��2(�?             6@������������������������       �                     4@������������������������       �                      @y       �                    �?�s�ۺ�?�             s@z       �       
             �?�>$�*��?            �D@{       �                    �?���Q��?             >@|       �                   �a@��
ц��?             :@}       ~                   @[@�G�z��?
             4@������������������������       �                     �?       �                   �a@D�n�3�?	             3@�       �                    �I@8�Z$���?             *@�       �                   @_@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    @H@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     &@�       �       	          ����?���:�?�            pp@�       �       
             �?P̏����?$            �L@�       �       	          ����?�ʈD��?            �E@������������������������       �                     @@�       �                    �?���|���?             &@�       �                   `]@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �\@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   `d@����X�?
             ,@�       �                   `c@X�<ݚ�?             "@�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?X�?٥�?�            �i@�       �                   �U@ �h�7W�?`            �c@������������������������       �                     �?�       �       
             �? �\���?_            �c@�       �                    �?��<�Ұ?W            `b@�       �                   Pb@@�n�1�?M            @_@�       �                    �? ��+&ɐ?J            @^@������������������������       �        5            �V@�       �                   �[@�g�y��?             ?@������������������������       �                     �?������������������������       �                     >@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �b@��2(&�?
             6@������������������������       �        	             3@������������������������       �                     @�       �                    �?���!pc�?             &@�       �                    @M@z�G�z�?             $@������������������������       �                     @�       �                    �N@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   @s@`Ql�R�?#            �G@������������������������       �                    �E@�       �                    �?      �?             @�       �       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�t�b�|D      h�h*h-K ��h/��R�(KK�KK��ha�B�       �t@     @y@     �q@     `b@      p@      Z@     �n@     @R@     �C@     �K@              6@     �C@     �@@      5@       @       @       @              �?       @      �?      @               @      �?       @                      �?      *@              2@      ?@      @      7@      @              @      7@      @      $@              "@      @      �?      @                      �?              *@      (@       @      &@       @      �?      �?      �?                      �?      $@      �?       @               @      �?              �?       @              �?      @      �?      �?              �?      �?                      @     �i@      2@     �i@      0@     �g@      (@      K@              a@      (@      @       @               @      @             �`@      $@     �`@      "@      E@       @      @      @              @      @              C@      @      "@      @      "@                      @      =@             �V@      �?     �L@              A@      �?      A@                      �?              �?      .@      @       @       @       @                       @      *@       @      (@              �?       @      �?                       @               @      &@      ?@      @      <@      @      @      @      �?      @              �?      �?              �?      �?                      @       @      8@              6@       @       @               @       @              @      @      @               @      @       @                      @      ;@     �E@      @      ?@      �?      9@      �?      �?      �?                      �?              8@      @      @      �?      @              @      �?      �?              �?      �?              @      �?              �?      @              6@      (@       @      $@              @       @      @              @       @              4@       @      4@                       @     �G@     p@      7@      2@      (@      2@      (@      ,@      &@      "@              �?      &@       @      &@       @      @       @      @                       @       @                      @      �?      @      �?                      @              @      &@              8@     �m@      ,@     �E@      @     �C@              @@      @      @      �?      @      �?                      @      @       @      @                       @      $@      @      @      @      @      �?              �?      @                      @      @              $@     �h@      "@     �b@      �?               @     �b@      @     �a@       @     �^@      �?      ^@             �V@      �?      >@      �?                      >@      �?      @      �?                      @      @      3@              3@      @              @       @       @       @              @       @      @       @                      @      �?              �?      G@             �E@      �?      @      �?       @      �?                       @              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�BHzhG        hNhG        hGKhHKhIh*h-K ��h/��R�(KK��ha�C              �?�t�bhUhfhPC       ���R�hjKhkhnKh*h-K ��h/��R�(KK��hP�C       �t�bK��R�}�(hKhxK�hyh*h-K ��h/��R�(KKŅ�h��B+         H       	          ����?�[��N�?�           ��@              
             �?��)��?�            �v@                          �_@��>4��?H             \@              	          hff�? pƵHP�?#             J@������������������������       �                    �G@                          �\@z�G�z�?             @������������������������       �                     @������������������������       �                     �?	                          pq@�z�G��?%             N@
              	          ����?�û��|�?             G@                           �?z�G�z�?             9@������������������������       �        	             .@                          �\@      �?             $@������������������������       �                      @                           �?      �?              @������������������������       �                     @                           �?      �?             @������������������������       �                     �?������������������������       �                     @                            O@�ՙ/�?             5@                           �?և���X�?	             ,@������������������������       �                     @                           �?�����H�?             "@������������������������       �                     @                           �?z�G�z�?             @              	            �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@        7                    �?0�|#�p�?�            �o@!       "                     B@R=6�z�?&            @P@������������������������       �                     @#       *                    T@r֛w���?$             O@$       )                   �\@d}h���?             ,@%       (                    �?      �?              @&       '                   �X@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @+       6       	          ����?8��8���?             H@,       5                    `@4?,R��?             B@-       4                   0e@�q�q�?             .@.       /                    �?r�q��?	             (@������������������������       �                     @0       3                    _@�<ݚ�?             "@1       2                   �g@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     5@������������������������       �                     (@8       E                    �Q@8�o+�?m            �g@9       D                   �g@�˫���?j             g@:       ;                    �?@i�)ԙ�?i            �f@������������������������       �                     �N@<       C                    �?��7�K¨?I            @^@=       @                   @[@�?�|�?B            �[@>       ?                   �_@����X�?             @������������������������       �                     @������������������������       �                      @A       B                   �t@�ջ����??             Z@������������������������       �        >            �Y@������������������������       �                     �?������������������������       �                     $@������������������������       �                      @F       G                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @I       �       
             �?ByL5���?�            �v@J       i                    �? ��om��?�            ps@K       `                    �?�q�q�?             E@L       _                     Q@�חF�P�?             ?@M       \                   �x@�r����?             >@N       [                    �? �Cc}�?             <@O       Z                   �`@R���Q�?             4@P       S                    _@      �?              @Q       R                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?T       U                    �I@�q�q�?             @������������������������       �                     @V       W                    �J@�q�q�?             @������������������������       �                     �?X       Y                    `@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             (@������������������������       �                      @]       ^                    �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?a       b                    �?"pc�
�?             &@������������������������       �                     @c       d       
             �?      �?              @������������������������       �                     �?e       h                   �b@����X�?             @f       g                    o@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?j       �                   �b@�E�J��?�            �p@k       �                    �?@�E~��?�            @o@l       �                   �z@�]��?�            �i@m       �                   Xp@XB���?�            `i@n       �                   �_@�U�e?Ƕ?]            �b@o       |                   �_@      �?=             X@p       w                    �?�>4և��?             <@q       r                   Ph@���}<S�?             7@������������������������       �                     0@s       v                     O@����X�?             @t       u       	             �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @x       {                    �?���Q��?             @y       z                    �O@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @}       ~                    �? ��ʻ��?,             Q@������������������������       �                     E@       �       	          ����? ��WV�?             :@�       �                   �`@z�G�z�?             @�       �                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     5@�       �                    \@@3����?              K@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     H@������������������������       �        #            �J@�       �                     L@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �`@��2(&�?             F@�       �                    c@(;L]n�?             >@������������������������       �                     8@�       �       	          hff @r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?X�Cc�?             ,@������������������������       �                     @�       �                     P@      �?             $@�       �                   �`@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    e@�����?             3@�       �                    `@�eP*L��?	             &@�       �                   Pl@r�q��?             @�       �       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �X@z�G�z�?             @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �B@      �?              @������������������������       �                     �?������������������������       �                     @�       �                   q@h�����?%             L@�       �                    _@\�Uo��?             C@������������������������       �                     $@�       �                    @N@���>4��?             <@�       �                    b@�û��|�?             7@�       �       	          033�?��.k���?             1@�       �                    �K@      �?              @������������������������       �                     @������������������������       �                      @�       �                    �?�<ݚ�?             "@�       �                    �?      �?              @������������������������       �                     @�       �                   @`@z�G�z�?             @�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   0b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�����H�?
             2@�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@�t�bh�h*h-K ��h/��R�(KK�KK��ha�BP       �s@     Pz@      o@     �]@      3@     @W@      �?     �I@             �G@      �?      @              @      �?              2@      E@      2@      <@      @      4@              .@      @      @               @      @      @      @              �?      @      �?                      @      *@       @      @       @      @              �?       @              @      �?      @      �?      @              @      �?                      �?      @                      ,@     �l@      :@      G@      3@              @      G@      0@      @      &@      @      @      @      @              @      @                      �?              @     �E@      @      ?@      @      $@      @      $@       @      @              @       @      @      �?              �?      @                      �?              @      5@              (@             �f@      @     `f@      @     `f@      @     �N@             �]@      @      [@      @      @       @      @                       @     �Y@      �?     �Y@                      �?      $@                       @      @       @      @                       @     @P@     �r@      A@     Pq@      ,@      <@      @      :@      @      :@      @      9@      @      1@      @      @      �?      �?              �?      �?               @      @              @       @      �?      �?              �?      �?              �?      �?                      (@               @      �?      �?              �?      �?              �?              "@       @      @              @       @      �?              @       @      @      �?      @                      �?              �?      4@      o@      ,@     �m@       @     �h@      @     �h@      @     �a@      @     �V@      @      7@       @      5@              0@       @      @       @       @       @                       @              @      @       @      �?       @      �?                       @       @              �?     �P@              E@      �?      9@      �?      @      �?      �?      �?                      �?              @              5@      �?     �J@      �?      @              @      �?                      H@             �J@      �?       @               @      �?              @      C@      �?      =@              8@      �?      @      �?                      @      @      "@              @      @      @      @      �?              �?      @                      @      @      *@      @      @      �?      @      �?       @               @      �?                      @      @      �?      �?      �?              �?      �?              @              �?      @      �?                      @      ?@      9@      .@      7@              $@      .@      *@      ,@      "@       @      "@      @       @      @                       @       @      @      �?      @              @      �?      @      �?      �?              �?      �?                      @      �?              @              �?      @              @      �?              0@       @      �?       @      �?                       @      .@        �t�bubhhubehhub.